magic
tech scmos
timestamp 1480861270
<< nwell >>
rect 1074 40 1078 45
rect 618 -142 626 -133
<< pwell >>
rect 729 317 739 321
<< metal1 >>
rect 194 1191 202 1199
rect 1074 1194 1082 1200
rect 1000 1168 1055 1180
rect 1000 1073 1055 1085
rect 1001 926 1056 938
rect 1230 924 1234 926
rect 200 892 208 898
rect 1000 881 1008 924
rect 1073 892 1078 899
rect 1872 881 1880 927
rect 1000 836 1055 848
rect 1001 748 1056 760
rect 201 590 208 596
rect 1001 581 1009 624
rect 1074 591 1083 597
rect 1871 580 1879 626
rect 1001 559 1056 571
rect 1001 480 1056 492
rect -35 456 -31 458
rect -35 453 -29 456
rect -33 366 -29 453
rect 1000 390 1055 402
rect -35 336 -31 339
rect -35 335 -29 336
rect -33 246 -29 335
rect 663 312 672 317
rect 200 290 207 296
rect 1000 279 1008 322
rect 1131 313 1132 319
rect 1127 308 1132 313
rect 1075 290 1087 298
rect 1872 278 1880 318
rect -35 217 -32 221
rect -35 134 -31 217
rect 1000 194 1055 206
rect 1000 128 1055 140
rect -34 120 -30 124
rect -34 97 -27 101
rect -33 57 -25 65
rect -33 17 -25 24
rect 999 23 1054 35
rect -33 16 -17 17
rect 311 16 331 22
rect -25 -6 -17 16
rect 13 -7 20 -3
rect 31 -7 39 -4
rect 42 -6 50 16
rect 80 -6 87 -3
rect 147 -8 154 -3
rect 176 -6 184 -5
rect 214 -10 221 -5
rect 244 -8 252 -5
rect 256 -6 260 -2
rect 282 -3 288 4
rect 282 -5 289 -3
rect 311 -5 319 16
rect 358 14 363 19
rect 381 12 389 17
rect 367 6 389 12
rect 340 -3 345 2
rect 300 -6 308 -5
rect 349 -6 356 3
rect 367 -5 375 6
rect 416 -5 423 12
rect 461 11 466 16
rect 483 -5 490 4
rect 551 5 558 12
rect 551 -7 558 -2
rect 1018 9 1024 11
rect 1018 6 1096 9
rect 618 -6 625 3
rect 647 -6 655 -5
rect 685 -8 692 4
rect 752 -5 759 3
rect 820 -7 827 4
rect 887 -7 894 4
rect 954 -5 961 4
rect 1021 -8 1028 2
rect 1089 -5 1096 6
rect 1099 5 1107 21
rect 1188 7 1195 33
rect 1574 22 1590 27
rect 1664 23 1672 24
rect 1768 23 1784 25
rect 1790 23 1828 31
rect 1099 -2 1126 5
rect 1118 -6 1126 -2
rect 1156 -1 1195 7
rect 1223 5 1230 6
rect 1156 -6 1163 -1
rect 1223 -5 1230 -1
rect 1290 2 1293 7
rect 1290 -3 1298 2
rect 1358 6 1397 12
rect 1404 6 1405 12
rect 1574 11 1580 22
rect 1290 -7 1297 -3
rect 1358 -7 1365 6
rect 1425 -6 1432 0
rect 1492 0 1506 7
rect 1559 6 1580 11
rect 1589 10 1622 19
rect 1492 -6 1499 0
rect 1559 -7 1566 6
rect 1589 -9 1597 10
rect 1664 8 1673 23
rect 1716 10 1724 22
rect 1768 17 1787 23
rect 1644 2 1673 8
rect 1694 6 1701 8
rect 1644 1 1672 2
rect 1627 -6 1634 -2
rect 1645 -9 1652 1
rect 1715 3 1731 10
rect 1693 -7 1701 -2
rect 1723 -8 1731 3
rect 1761 -6 1768 -1
rect 1779 -7 1787 17
rect 1790 -7 1798 23
rect 1870 17 1922 24
rect 1896 4 1902 8
rect 1828 -5 1835 -2
rect 1896 -8 1902 -3
rect 1914 -6 1922 17
rect 2097 6 2104 12
rect 1963 -5 1970 -1
rect 2030 -5 2037 -2
rect 2097 -6 2104 0
<< m2contact >>
rect 1127 605 1132 610
rect 1127 302 1132 308
rect 31 57 39 65
rect 1188 33 1195 40
rect 31 -4 39 4
rect 214 -5 221 1
<< metal2 >>
rect 255 1188 259 1201
rect 461 1195 465 1201
rect 564 1195 568 1201
rect 667 1196 671 1201
rect 770 1196 774 1201
rect 873 1196 877 1201
rect 975 1198 980 1201
rect 358 1188 362 1192
rect 975 1160 978 1198
rect 979 1189 980 1197
rect 228 605 1127 610
rect 131 302 157 308
rect 169 88 175 326
rect 217 302 1127 308
rect 165 82 175 88
rect 31 4 39 57
rect 165 58 171 82
rect 165 52 175 58
rect 169 23 175 52
rect 214 41 1074 45
rect 214 40 848 41
rect 867 40 1074 41
rect 122 17 175 23
rect 122 12 128 17
rect 4 -5 9 1
rect 71 8 128 12
rect 71 -6 76 8
rect 138 -6 143 4
rect 205 -6 210 21
rect 214 1 221 40
rect 1195 39 1474 40
rect 1195 33 1473 39
rect 357 22 362 26
rect 357 16 456 22
rect 999 19 1030 28
rect 999 17 1007 19
rect 273 -6 278 2
rect 282 -3 288 4
rect 340 -6 345 2
rect 416 5 423 12
rect 407 -7 412 4
rect 451 2 456 16
rect 461 11 466 16
rect 451 -3 479 2
rect 483 -3 490 4
rect 474 -6 479 -3
rect 542 -8 547 3
rect 551 5 558 12
rect 781 8 791 17
rect 801 8 1007 17
rect 1023 14 1030 19
rect 1341 18 1421 22
rect 1023 7 1108 14
rect 1023 6 1054 7
rect 1099 6 1108 7
rect 1249 16 1421 18
rect 1249 12 1347 16
rect 609 -6 614 3
rect 618 -3 625 3
rect 685 -3 692 4
rect 752 -3 759 3
rect 676 -5 681 -3
rect 743 -5 748 -3
rect 811 -6 816 2
rect 820 -3 827 4
rect 878 -7 883 3
rect 887 -3 894 4
rect 945 -7 950 2
rect 954 -2 961 4
rect 1021 -3 1028 2
rect 1012 -7 1017 -3
rect 1080 -6 1085 3
rect 1099 -1 1143 6
rect 1138 -7 1152 -1
rect 1214 -6 1219 6
rect 1223 5 1230 6
rect 1263 -1 1287 7
rect 1281 -6 1287 -1
rect 1349 -1 1363 5
rect 1349 -6 1354 -1
rect 1416 -7 1421 16
rect 1476 -2 1488 5
rect 1483 -6 1488 -2
rect 1550 -6 1555 -1
rect 1618 -7 1623 5
rect 1685 -7 1690 -1
rect 1752 -6 1757 -2
rect 1819 -5 1824 -3
rect 1887 -6 1892 -2
rect 1954 -5 1959 5
rect 2021 -6 2026 4
rect 2092 1 2093 11
rect 2087 -5 2093 1
rect 90 -242 95 -238
rect 359 -242 364 -238
rect 628 -242 633 -237
rect 897 -242 902 -235
rect 1166 -247 1171 -234
rect 1435 -246 1440 -235
rect 1704 -247 1710 -236
rect 1973 -242 1978 -235
<< m3contact >>
rect 222 605 228 610
rect 124 302 131 308
rect 157 302 164 308
rect 175 321 181 326
rect 210 302 217 308
rect 4 1 9 6
rect 1074 40 1079 45
rect 204 21 210 27
rect 138 4 143 9
rect 1473 32 1481 39
rect 268 -3 273 2
rect 335 -3 340 2
rect 407 4 412 10
rect 542 3 547 9
rect 791 8 801 17
rect 604 -3 609 3
rect 806 -3 811 2
rect 873 -3 878 3
rect 940 -3 945 2
rect 1075 -3 1080 3
rect 1254 -1 1263 8
rect 1363 -1 1368 5
rect 1467 -2 1476 5
rect 1550 -1 1555 4
rect 1613 0 1618 5
rect 1685 -1 1690 5
rect 1748 -2 1757 5
rect 1819 -3 1824 2
rect 1887 -2 1892 3
rect 2014 -3 2021 4
rect 2083 1 2092 11
rect 582 -175 587 -170
<< m123contact >>
rect -14 365 -8 370
rect -26 246 -20 251
rect -36 128 -30 134
rect 658 312 663 317
rect 13 -3 20 4
rect 80 -3 87 4
rect 147 -3 154 3
rect 1590 22 1595 27
rect 288 -3 295 4
rect 356 -2 363 5
rect 423 5 430 12
rect 461 6 466 11
rect 483 4 490 11
rect 551 -2 558 5
rect 618 3 625 10
rect 1012 6 1018 11
rect 676 -3 681 2
rect 692 -3 699 4
rect 827 -3 834 4
rect 894 -3 901 4
rect 961 -2 968 4
rect 1028 -3 1035 2
rect 1223 -1 1230 5
rect 1293 2 1298 7
rect 1397 6 1404 12
rect 1425 0 1432 7
rect 1506 0 1514 7
rect 1627 -2 1634 5
rect 1694 -2 1703 6
rect 1761 -1 1768 6
rect 1828 -2 1835 3
rect 1896 -3 1902 4
rect 1963 -1 1970 5
rect 2030 -2 2037 4
rect 2097 0 2104 6
rect 53 -175 58 -170
rect 322 -175 327 -170
rect 591 -175 596 -170
rect 860 -175 865 -170
rect 1129 -175 1134 -170
rect 1398 -175 1403 -170
rect 1667 -175 1672 -170
rect 1936 -175 1941 -170
<< metal3 >>
rect 131 924 212 929
rect 131 501 137 924
rect 4 495 137 501
rect 141 907 245 915
rect 616 907 656 915
rect 141 809 149 907
rect -36 3 -30 128
rect -26 17 -20 246
rect -14 -7 -8 365
rect 4 6 9 495
rect 141 491 148 809
rect 13 485 148 491
rect 152 623 213 628
rect 13 4 20 485
rect 152 481 157 623
rect 138 475 157 481
rect 163 605 222 610
rect 80 302 124 308
rect 80 4 87 302
rect 138 9 143 475
rect 163 471 169 605
rect 147 466 169 471
rect 147 3 153 466
rect 181 321 213 326
rect 588 319 596 534
rect 164 302 210 308
rect 1012 11 1018 891
rect -14 -8 2088 -7
rect -13 -12 2088 -8
rect -36 -170 -30 -28
rect 32 -29 2123 -23
rect -24 -43 2066 -37
rect -26 -102 -20 -61
rect -26 -107 2008 -102
rect -36 -175 53 -170
rect 58 -175 322 -170
rect 327 -175 582 -170
rect 587 -175 591 -170
rect 596 -175 860 -170
rect 865 -175 1129 -170
rect 1134 -175 1398 -170
rect 1403 -175 1667 -170
rect 1672 -175 1936 -170
<< m234contact >>
rect 1209 6 1219 13
rect 1242 12 1249 18
rect 743 -3 748 2
rect 1012 -3 1017 2
rect 1946 -3 1954 5
<< m4contact >>
rect 622 922 630 929
rect 720 924 728 930
rect 821 924 831 932
rect 1076 924 1084 933
rect 1488 924 1495 932
rect 245 907 254 915
rect 606 907 616 915
rect 656 907 666 915
rect -26 11 -20 17
rect -36 -3 -30 3
rect 308 623 315 629
rect 588 534 596 541
rect 529 20 536 26
rect 627 20 633 26
rect 835 23 847 35
rect 461 11 466 16
rect 1718 621 1726 629
rect 1594 322 1602 327
rect 1710 22 1716 28
rect 1425 7 1432 14
rect 1828 3 1835 8
rect 1805 -3 1819 2
rect 2072 1 2083 11
rect 2097 6 2104 12
rect -36 -28 -30 -22
rect -26 -61 -20 -55
<< metal4 >>
rect 236 954 729 962
rect 720 930 729 954
rect 728 926 729 930
rect 821 932 831 995
rect 254 907 606 915
rect 622 903 630 922
rect 661 915 741 916
rect 1076 915 1084 924
rect 666 907 1084 915
rect 1488 909 1494 924
rect 401 897 630 903
rect 1291 902 1494 909
rect 925 676 935 705
rect 1209 691 1741 694
rect 1209 683 1730 691
rect 1181 642 1888 650
rect 308 613 315 623
rect 268 607 315 613
rect 424 610 456 611
rect 471 610 1067 611
rect 424 605 1067 610
rect 1718 604 1726 621
rect 634 596 662 601
rect 1718 595 1761 604
rect 1876 592 1888 642
rect 529 590 586 591
rect 536 583 586 590
rect 579 541 586 583
rect 1876 582 1889 592
rect 579 534 588 541
rect 1170 451 1397 452
rect 1615 451 1787 452
rect 1170 443 1787 451
rect 1170 441 1795 443
rect 1390 440 1627 441
rect 1175 350 1684 357
rect 356 302 991 308
rect 1296 301 1453 311
rect 1594 219 1602 322
rect 1425 212 1602 219
rect 1425 124 1432 212
rect 1425 117 1441 124
rect 1081 87 1421 88
rect 993 86 1421 87
rect 735 81 1421 86
rect 735 80 1133 81
rect 735 79 1039 80
rect 461 65 748 70
rect 1434 68 1441 117
rect 1876 116 1890 582
rect 1454 82 1547 88
rect 1454 81 1555 82
rect 461 16 466 65
rect -36 -22 -30 -3
rect -26 -55 -20 11
rect 288 -3 289 4
rect 269 -29 406 -22
rect 529 -34 536 20
rect 627 14 633 20
rect 627 9 725 14
rect 718 5 725 9
rect 743 2 748 65
rect 1424 62 1441 68
rect 1877 62 1890 116
rect 764 41 1249 48
rect 764 40 848 41
rect 867 40 1249 41
rect 847 23 857 35
rect 1242 18 1249 40
rect 814 17 1010 18
rect 814 14 1017 17
rect 814 13 1099 14
rect 814 9 1209 13
rect 811 8 1209 9
rect 967 7 1209 8
rect 1091 6 1209 7
rect 1425 14 1432 62
rect 1877 59 2008 62
rect 1878 49 2008 59
rect 1795 37 2104 41
rect 1795 34 1796 37
rect 1803 34 2104 37
rect 1716 22 1836 28
rect 1828 8 1835 22
rect 2097 12 2104 34
rect 1828 -1 1835 3
rect 1929 -3 1946 5
rect 2072 -3 2083 1
rect 572 -20 876 -14
rect 587 -29 943 -24
rect 1012 -34 1017 -3
rect 529 -40 1017 -34
rect 529 -41 536 -40
rect 1080 -45 1085 -3
rect 402 -50 1085 -45
rect 726 -69 1263 -60
rect 255 -91 539 -82
rect 1125 -83 1348 -82
rect 255 -92 442 -91
rect 962 -91 1348 -83
rect 962 -92 1138 -91
rect 895 -104 1322 -96
rect 1146 -109 1302 -108
rect 828 -116 1302 -109
rect 759 -127 1280 -120
rect 1302 -127 1491 -120
rect 626 -141 1162 -133
rect 618 -142 1162 -141
rect 490 -156 1175 -148
rect 1376 -160 1382 -159
rect 1028 -168 1382 -160
rect 692 -179 1146 -173
rect 684 -180 1146 -179
rect 1156 -180 1159 -173
rect 238 -193 1368 -186
rect 845 -207 1456 -200
rect 835 -208 1456 -207
rect 1805 -214 1818 -3
rect 1336 -215 1569 -214
rect 1793 -215 1818 -214
rect 1104 -216 1818 -215
rect 871 -226 1818 -216
rect 1929 -222 1939 -3
rect 2072 -13 2082 -3
rect 1945 -25 2082 -13
rect 1945 -26 2079 -25
rect 871 -227 1337 -226
rect 1562 -227 1795 -226
rect 871 -228 1104 -227
rect 1929 -232 1938 -222
rect 1197 -233 1663 -232
rect 1871 -233 1938 -232
rect 980 -244 1938 -233
rect 968 -245 1201 -244
rect 1659 -245 1938 -244
rect 932 -251 1439 -250
rect 1945 -251 1958 -26
rect 932 -258 1958 -251
rect 1422 -259 1958 -258
<< m345contact >>
rect 411 935 416 944
rect 308 924 314 930
rect 526 923 534 930
rect 1590 938 1600 948
rect 926 925 936 933
rect 1179 925 1186 931
rect 1282 925 1290 931
rect 1384 924 1393 934
rect 1695 924 1702 930
rect 1801 924 1816 934
rect 1012 891 1018 900
rect 437 623 442 628
rect 529 622 536 629
rect 627 623 634 628
rect 733 623 741 629
rect 842 624 855 633
rect 949 623 958 629
rect 1194 623 1202 630
rect 1282 624 1290 632
rect 1404 618 1414 629
rect 1489 624 1501 636
rect 1588 627 1597 635
rect 1820 623 1829 630
rect 340 320 345 325
rect 437 319 443 324
rect 538 316 546 323
rect 588 312 596 319
rect 729 317 739 325
rect 844 320 853 325
rect 939 319 948 325
rect 1179 322 1186 328
rect 1282 322 1293 330
rect 1384 322 1400 334
rect 1486 324 1496 333
rect 653 312 658 317
rect 1694 321 1704 329
rect 1821 322 1829 329
rect 416 5 423 12
rect 273 -3 278 2
rect 282 -3 288 4
rect 340 -3 345 2
rect 349 -2 356 4
rect 407 -2 412 4
rect 483 -3 491 4
rect 728 21 735 28
rect 551 5 558 12
rect 542 -3 547 3
rect 609 -3 614 3
rect 618 -3 625 3
rect 671 -3 676 2
rect 685 -3 692 4
rect 935 22 945 29
rect 1175 22 1184 31
rect 781 8 791 17
rect 1280 22 1289 29
rect 1384 22 1395 30
rect 1473 39 1481 46
rect 1796 32 1803 37
rect 1491 21 1501 28
rect 1223 5 1230 12
rect 752 -3 759 3
rect 811 -3 816 2
rect 820 -3 827 4
rect 878 -3 883 3
rect 887 -3 894 4
rect 945 -3 950 2
rect 954 -2 961 4
rect 1021 -3 1028 2
rect 1080 -3 1085 3
rect 1263 -1 1272 8
rect 1404 6 1411 12
rect 1293 -3 1298 2
rect 1368 -1 1374 5
rect 1458 -2 1467 5
rect 1514 0 1522 7
rect 1550 4 1555 9
rect 1627 5 1634 12
rect 1685 5 1690 11
rect 1694 6 1703 14
rect 1761 6 1768 13
rect 1607 0 1613 5
rect 1740 -2 1748 5
rect 1896 4 1902 11
rect 1963 5 1970 11
rect 1882 -2 1887 3
rect 2014 4 2021 11
rect 2030 4 2037 10
<< m5contact >>
rect 821 995 831 1005
rect 223 951 236 966
rect 393 896 401 903
rect 1283 902 1291 909
rect 923 705 936 719
rect 1188 682 1209 696
rect 1730 681 1742 691
rect 922 662 935 676
rect 1171 633 1181 650
rect 262 607 268 613
rect 416 605 424 611
rect 1067 605 1074 611
rect 627 596 634 601
rect 662 596 670 601
rect 1761 595 1768 604
rect 529 583 536 590
rect 1152 441 1170 453
rect 1787 443 1798 453
rect 1168 349 1175 357
rect 1684 350 1690 357
rect 349 302 356 308
rect 991 302 997 308
rect 1283 300 1296 311
rect 1453 301 1465 311
rect 728 79 735 86
rect 1421 81 1429 88
rect 1446 81 1454 88
rect 1547 82 1555 89
rect 262 -29 269 -22
rect 406 -29 413 -22
rect 718 -1 725 5
rect 752 39 764 48
rect 857 23 869 35
rect 804 9 814 19
rect 2008 49 2021 62
rect 565 -20 572 -14
rect 876 -20 883 -14
rect 579 -29 587 -24
rect 943 -29 950 -23
rect 394 -51 402 -44
rect 718 -69 726 -60
rect 1263 -69 1272 -60
rect 245 -92 255 -81
rect 539 -91 547 -82
rect 954 -92 962 -83
rect 1348 -91 1359 -82
rect 887 -104 895 -96
rect 1322 -104 1335 -96
rect 820 -116 828 -108
rect 1302 -116 1311 -108
rect 752 -127 759 -120
rect 1280 -127 1289 -120
rect 1293 -127 1302 -120
rect 1491 -127 1501 -120
rect 618 -141 626 -132
rect 1162 -142 1171 -133
rect 482 -156 490 -147
rect 1175 -156 1184 -146
rect 1020 -168 1028 -160
rect 1382 -168 1395 -158
rect 682 -179 692 -171
rect 1146 -180 1156 -172
rect 223 -195 238 -183
rect 1368 -193 1374 -186
rect 834 -207 845 -197
rect 1456 -208 1468 -200
rect 859 -228 871 -215
rect 968 -244 980 -232
rect 922 -258 932 -247
<< metal5 >>
rect 831 996 1616 1005
rect 427 989 435 990
rect 427 980 1187 989
rect 226 832 235 951
rect 245 935 411 944
rect 226 -183 236 832
rect 245 -81 255 935
rect 273 924 308 930
rect 262 -22 268 607
rect 273 2 278 924
rect 427 915 435 980
rect 282 907 435 915
rect 440 970 1165 976
rect 282 4 289 907
rect 440 903 447 970
rect 925 933 936 934
rect 394 868 401 896
rect 428 898 447 903
rect 526 907 534 923
rect 925 925 926 933
rect 526 899 648 907
rect 288 -3 289 4
rect 340 2 345 320
rect 349 4 356 302
rect 394 -44 402 868
rect 416 510 424 605
rect 416 12 423 510
rect 428 477 433 898
rect 437 618 442 623
rect 437 613 466 618
rect 461 559 466 613
rect 529 590 536 622
rect 627 601 634 623
rect 461 551 636 559
rect 427 466 433 477
rect 427 263 432 466
rect 437 331 616 338
rect 437 324 443 331
rect 538 323 546 326
rect 538 315 546 316
rect 538 308 574 315
rect 427 54 434 263
rect 565 245 574 308
rect 579 312 588 319
rect 427 47 558 54
rect 551 12 558 47
rect 407 -22 412 -2
rect 482 -78 491 -3
rect 482 -147 490 -78
rect 542 -82 547 -3
rect 565 -14 573 245
rect 572 -20 573 -14
rect 579 -24 587 312
rect 609 285 614 331
rect 608 271 614 285
rect 608 100 613 271
rect 608 97 614 100
rect 609 3 614 97
rect 630 2 636 551
rect 640 14 647 899
rect 925 719 936 925
rect 1158 921 1165 970
rect 1178 931 1187 980
rect 1424 939 1590 946
rect 1178 927 1179 931
rect 1186 927 1187 931
rect 1282 921 1290 925
rect 1158 913 1290 921
rect 1303 924 1384 934
rect 1012 902 1283 909
rect 1012 900 1018 902
rect 842 695 855 696
rect 842 684 1188 695
rect 842 633 855 684
rect 732 623 733 629
rect 924 646 935 662
rect 662 369 670 596
rect 732 389 741 623
rect 924 463 936 646
rect 949 643 957 644
rect 948 635 1171 643
rect 949 629 957 635
rect 1067 633 1171 635
rect 1194 611 1202 623
rect 1074 605 1202 611
rect 1212 624 1282 632
rect 1212 600 1221 624
rect 925 451 936 463
rect 1190 592 1221 600
rect 925 441 1152 451
rect 925 440 1162 441
rect 732 379 836 389
rect 827 374 836 379
rect 662 357 814 369
rect 653 337 790 343
rect 653 317 658 337
rect 739 320 763 321
rect 739 317 764 320
rect 729 314 764 317
rect 753 280 764 314
rect 780 297 790 337
rect 728 28 735 79
rect 752 48 764 280
rect 781 17 790 297
rect 804 19 814 357
rect 827 34 837 374
rect 844 357 854 358
rect 844 349 1168 357
rect 844 325 854 349
rect 853 320 854 325
rect 937 325 977 329
rect 937 320 939 325
rect 948 320 977 325
rect 827 32 845 34
rect 827 23 846 32
rect 640 9 768 14
rect 630 -3 671 2
rect 618 -132 625 -3
rect 685 -112 692 -3
rect 718 -60 725 -1
rect 763 2 768 9
rect 763 -3 811 2
rect 684 -171 692 -112
rect 752 -120 759 -3
rect 820 -108 827 -3
rect 835 -197 845 23
rect 857 10 869 23
rect 835 -209 845 -207
rect 858 -131 869 10
rect 922 29 939 30
rect 922 22 935 29
rect 878 -14 883 -3
rect 887 -96 894 -3
rect 858 -215 870 -131
rect 922 -247 932 22
rect 945 -23 950 -3
rect 954 -83 961 -2
rect 968 -232 977 320
rect 1136 322 1179 328
rect 1136 308 1143 322
rect 1190 309 1198 592
rect 1303 516 1312 924
rect 1302 510 1312 516
rect 1404 569 1414 618
rect 997 302 1143 308
rect 1147 302 1198 309
rect 1203 322 1282 330
rect 1021 -116 1028 -3
rect 1147 -112 1156 302
rect 1203 298 1211 322
rect 1162 289 1211 298
rect 1224 302 1283 311
rect 1021 -146 1029 -116
rect 1021 -160 1028 -146
rect 1146 -172 1157 -112
rect 1162 -133 1171 289
rect 1224 183 1231 302
rect 1223 176 1231 183
rect 1175 -146 1184 22
rect 1223 12 1230 176
rect 1263 -60 1272 -1
rect 1280 -120 1289 22
rect 1293 2 1298 5
rect 1293 -120 1298 -3
rect 1302 -108 1311 510
rect 1404 441 1413 569
rect 1404 435 1414 441
rect 1322 334 1335 336
rect 1321 322 1384 334
rect 1322 -96 1335 322
rect 1405 314 1414 435
rect 1346 304 1414 314
rect 1346 135 1359 304
rect 1404 236 1411 237
rect 1424 236 1434 939
rect 1453 636 1464 641
rect 1452 624 1489 636
rect 1501 624 1503 636
rect 1586 633 1588 634
rect 1513 627 1588 633
rect 1513 626 1595 627
rect 1513 625 1588 626
rect 1453 612 1464 624
rect 1453 311 1463 612
rect 1474 324 1486 332
rect 1474 323 1496 324
rect 1453 300 1463 301
rect 1404 228 1439 236
rect 1404 177 1411 228
rect 1424 226 1434 228
rect 1404 176 1412 177
rect 1347 -55 1359 135
rect 1405 67 1412 176
rect 1429 81 1446 88
rect 1454 81 1455 88
rect 1404 61 1412 67
rect 1348 -82 1359 -55
rect 1156 -180 1157 -172
rect 1368 -186 1374 -1
rect 1385 -158 1395 22
rect 1404 12 1411 61
rect 1474 46 1482 323
rect 1481 39 1482 46
rect 1474 33 1482 39
rect 1458 -200 1467 -2
rect 1491 -120 1501 21
rect 1515 7 1522 625
rect 1550 9 1555 82
rect 1607 5 1613 996
rect 1625 924 1695 930
rect 1626 922 1701 924
rect 1627 12 1634 922
rect 1733 691 1741 694
rect 1733 603 1741 681
rect 1684 11 1690 350
rect 1684 8 1685 11
rect 1694 14 1703 321
rect 1732 307 1741 603
rect 1731 296 1741 307
rect 1731 0 1740 296
rect 1761 13 1768 595
rect 1788 49 1797 443
rect 1803 377 1815 924
rect 1820 583 1829 623
rect 1820 572 1851 583
rect 1802 375 1815 377
rect 1802 67 1814 375
rect 1822 329 1832 330
rect 1829 322 1832 329
rect 1821 79 1832 322
rect 1840 91 1851 572
rect 1840 83 2038 91
rect 1821 71 1971 79
rect 1802 66 1869 67
rect 1802 65 1876 66
rect 1802 57 1878 65
rect 1813 56 1878 57
rect 1859 49 1867 51
rect 1787 41 1867 49
rect 1732 -2 1740 0
rect 1859 3 1867 41
rect 1871 17 1878 56
rect 1871 11 1902 17
rect 1963 11 1970 71
rect 2014 11 2021 49
rect 2030 10 2038 83
rect 2037 8 2038 10
rect 1859 -2 1882 3
rect 1887 -2 1891 3
rect 1458 -209 1467 -208
use decoder_and_memory  decoder_and_memory_0
timestamp 1480861270
transform 1 0 -65 0 1 14
box 30 -10 1945 1187
use mux81  mux81_0
timestamp 1480738159
transform 0 1 175 -1 0 -5
box 0 -204 237 65
use mux81  mux81_1
timestamp 1480738159
transform 0 1 444 -1 0 -5
box 0 -204 237 65
use mux81  mux81_2
timestamp 1480738159
transform 0 1 713 -1 0 -5
box 0 -204 237 65
use mux81  mux81_3
timestamp 1480738159
transform 0 1 982 -1 0 -5
box 0 -204 237 65
use mux81  mux81_4
timestamp 1480738159
transform 0 1 1251 -1 0 -5
box 0 -204 237 65
use mux81  mux81_5
timestamp 1480738159
transform 0 1 1520 -1 0 -5
box 0 -204 237 65
use mux81  mux81_6
timestamp 1480738159
transform 0 1 1789 -1 0 -5
box 0 -204 237 65
use mux81  mux81_7
timestamp 1480738159
transform 0 1 2058 -1 0 -5
box 0 -204 237 65
<< labels >>
rlabel metal1 -31 61 -31 61 3 Vdd
rlabel metal1 -31 19 -31 19 3 Gnd
rlabel metal2 92 -241 92 -241 1 out7
rlabel metal2 257 1191 257 1191 1 new7
rlabel metal2 360 1190 360 1190 1 new6
rlabel metal1 197 1196 197 1196 5 clk0
rlabel metal1 1076 1197 1076 1197 5 clk4
rlabel metal1 202 894 202 894 1 clk1
rlabel metal1 205 592 205 592 1 clk2
rlabel metal1 202 293 202 293 1 clk3
rlabel metal1 1076 296 1076 296 1 clk7
rlabel metal1 1076 596 1076 596 1 clk6
rlabel metal1 1074 898 1074 898 1 clk5
rlabel metal1 -34 456 -34 456 3 input2_r
rlabel metal1 -34 337 -34 337 3 input1_r
rlabel metal1 -34 219 -34 219 3 input0_r
rlabel metal1 -33 122 -33 122 3 clear_r
rlabel metal1 -33 99 -33 99 3 calc_hist_r
rlabel metal2 361 -241 361 -241 1 out6
rlabel metal2 630 -241 630 -241 1 out5
rlabel metal2 899 -240 899 -240 1 out4
rlabel metal2 1168 -246 1168 -246 1 out3
rlabel metal2 1437 -245 1437 -245 1 out2
rlabel metal2 1707 -246 1707 -246 1 out1
rlabel metal2 1973 -242 1978 -235 1 out0
rlabel metal2 978 1200 978 1200 5 new0
rlabel metal2 874 1200 874 1200 5 new1
rlabel metal2 770 1196 774 1201 5 new2
rlabel metal2 668 1200 668 1200 5 new3
rlabel metal2 565 1200 565 1200 5 new4
rlabel metal2 462 1200 462 1200 5 new5
<< end >>
