magic
tech scmos
timestamp 1480480681
<< nwell >>
rect -36 -3 140 28
rect -36 -84 140 -52
<< pwell >>
rect -36 -52 140 -3
<< ntransistor >>
rect -23 -13 -21 -9
rect 28 -13 30 -9
rect 70 -13 72 -9
rect 88 -13 90 -9
rect 104 -13 106 -9
rect 125 -13 127 -9
rect -25 -46 -23 -42
rect -5 -46 -3 -42
rect 23 -46 25 -42
rect 34 -46 36 -42
rect 81 -46 83 -42
rect 91 -46 93 -42
rect 108 -46 110 -42
<< ptransistor >>
rect -23 3 -21 9
rect 28 3 30 9
rect 70 3 72 9
rect 88 3 90 9
rect 104 3 106 9
rect 125 3 127 9
rect -25 -64 -23 -58
rect -5 -64 -3 -58
rect 23 -64 25 -58
rect 34 -64 36 -58
rect 81 -64 83 -58
rect 91 -64 93 -58
rect 108 -64 110 -58
<< ndiffusion >>
rect -24 -13 -23 -9
rect -21 -13 -19 -9
rect 27 -13 28 -9
rect 30 -13 33 -9
rect 69 -13 70 -9
rect 72 -13 75 -9
rect 87 -13 88 -9
rect 90 -13 91 -9
rect 103 -13 104 -9
rect 106 -13 109 -9
rect 124 -13 125 -9
rect 127 -13 130 -9
rect -26 -46 -25 -42
rect -23 -46 -20 -42
rect -6 -46 -5 -42
rect -3 -46 0 -42
rect 22 -46 23 -42
rect 25 -46 26 -42
rect 30 -46 34 -42
rect 36 -46 41 -42
rect 80 -46 81 -42
rect 83 -46 84 -42
rect 88 -46 91 -42
rect 93 -46 94 -42
rect 106 -46 108 -42
rect 110 -46 113 -42
<< pdiffusion >>
rect -28 8 -23 9
rect -24 4 -23 8
rect -28 3 -23 4
rect -21 8 -15 9
rect -21 4 -19 8
rect -21 3 -15 4
rect 23 8 28 9
rect 27 4 28 8
rect 23 3 28 4
rect 30 8 37 9
rect 30 4 33 8
rect 30 3 37 4
rect 65 8 70 9
rect 69 4 70 8
rect 65 3 70 4
rect 72 8 79 9
rect 72 4 75 8
rect 72 3 79 4
rect 83 8 88 9
rect 87 4 88 8
rect 83 3 88 4
rect 90 8 95 9
rect 90 4 91 8
rect 90 3 95 4
rect 99 8 104 9
rect 103 4 104 8
rect 99 3 104 4
rect 106 8 113 9
rect 106 4 109 8
rect 106 3 113 4
rect 120 8 125 9
rect 124 4 125 8
rect 120 3 125 4
rect 127 8 134 9
rect 127 4 130 8
rect 127 3 134 4
rect -30 -59 -25 -58
rect -26 -63 -25 -59
rect -30 -64 -25 -63
rect -23 -59 -16 -58
rect -23 -63 -20 -59
rect -23 -64 -16 -63
rect -10 -59 -5 -58
rect -6 -63 -5 -59
rect -10 -64 -5 -63
rect -3 -59 4 -58
rect -3 -63 0 -59
rect -3 -64 4 -63
rect 22 -64 23 -58
rect 25 -64 26 -58
rect 30 -64 34 -58
rect 36 -64 41 -58
rect 80 -64 81 -58
rect 83 -64 84 -58
rect 88 -64 91 -58
rect 93 -64 94 -58
rect 106 -64 108 -58
rect 110 -64 113 -58
<< ndcontact >>
rect -28 -13 -24 -9
rect -19 -13 -15 -9
rect 23 -13 27 -9
rect 33 -13 37 -9
rect 65 -13 69 -9
rect 75 -13 79 -9
rect 83 -13 87 -9
rect 91 -13 95 -9
rect 99 -13 103 -9
rect 109 -13 113 -9
rect 120 -13 124 -9
rect 130 -13 134 -9
rect -30 -46 -26 -42
rect -20 -46 -16 -42
rect -10 -46 -6 -42
rect 0 -46 4 -42
rect 18 -46 22 -42
rect 26 -46 30 -42
rect 41 -46 45 -42
rect 76 -46 80 -42
rect 84 -46 88 -42
rect 94 -46 98 -42
rect 102 -46 106 -42
rect 113 -46 117 -42
<< pdcontact >>
rect -28 4 -24 8
rect -19 4 -15 8
rect 23 4 27 8
rect 33 4 37 8
rect 65 4 69 8
rect 75 4 79 8
rect 83 4 87 8
rect 91 4 95 8
rect 99 4 103 8
rect 109 4 113 8
rect 120 4 124 8
rect 130 4 134 8
rect -30 -63 -26 -59
rect -20 -63 -16 -59
rect -10 -63 -6 -59
rect 0 -63 4 -59
rect 18 -64 22 -58
rect 26 -64 30 -58
rect 41 -64 45 -58
rect 76 -64 80 -58
rect 84 -64 88 -58
rect 94 -64 98 -58
rect 102 -64 106 -58
rect 113 -64 117 -58
<< psubstratepcontact >>
rect -24 -29 -20 -25
rect 35 -29 39 -25
rect 92 -29 96 -25
rect 125 -29 129 -25
<< nsubstratencontact >>
rect 7 21 11 25
rect 80 21 84 25
rect 120 21 124 25
rect 7 -81 11 -77
rect 60 -81 64 -77
rect 98 -81 102 -77
<< polysilicon >>
rect -23 9 -21 12
rect 28 9 30 12
rect 70 9 72 12
rect 88 9 90 12
rect 104 9 106 12
rect 125 9 127 12
rect -23 0 -21 3
rect 28 -1 30 3
rect 70 -1 72 3
rect 88 0 90 3
rect 104 -1 106 3
rect 125 -1 127 3
rect -23 -9 -21 -6
rect 28 -9 30 -5
rect 70 -9 72 -5
rect 88 -9 90 -6
rect 104 -9 106 -5
rect 125 -9 127 -5
rect -23 -16 -21 -13
rect 28 -16 30 -13
rect 70 -16 72 -13
rect 88 -16 90 -13
rect 104 -16 106 -13
rect 125 -16 127 -13
rect -25 -42 -23 -39
rect -5 -42 -3 -39
rect 23 -42 25 -38
rect 34 -42 36 -39
rect 81 -42 83 -38
rect 91 -42 93 -39
rect 108 -42 110 -39
rect -25 -51 -23 -46
rect -5 -51 -3 -46
rect 23 -49 25 -46
rect 34 -51 36 -46
rect 81 -49 83 -46
rect 91 -51 93 -46
rect 108 -51 110 -46
rect -25 -58 -23 -55
rect -5 -58 -3 -55
rect 23 -58 25 -55
rect 34 -58 36 -55
rect 81 -58 83 -55
rect 91 -58 93 -55
rect 108 -58 110 -55
rect -25 -67 -23 -64
rect -5 -67 -3 -64
rect 23 -68 25 -64
rect 34 -67 36 -64
rect 81 -68 83 -64
rect 91 -67 93 -64
rect 108 -67 110 -64
<< polycontact >>
rect -23 12 -19 16
rect 86 12 90 16
rect 26 -5 30 -1
rect 68 -5 72 -1
rect 102 -5 106 -1
rect 123 -5 127 -1
rect -23 -20 -19 -16
rect 86 -20 90 -16
rect 21 -38 25 -34
rect 79 -38 83 -34
rect -27 -55 -23 -51
rect -7 -55 -3 -51
rect 34 -55 38 -51
rect 91 -55 95 -51
rect 106 -55 110 -51
rect 21 -72 25 -68
rect 79 -72 83 -68
<< metal1 >>
rect -30 25 127 27
rect -30 21 7 25
rect 11 21 80 25
rect 84 21 120 25
rect 124 21 127 25
rect -30 20 127 21
rect -30 19 76 20
rect 87 19 127 20
rect -19 12 -3 16
rect -28 8 -24 9
rect -28 1 -24 4
rect -36 -3 -24 1
rect -28 -9 -24 -3
rect -19 8 -15 9
rect -19 -1 -15 4
rect 23 8 27 19
rect 23 3 27 4
rect 33 8 37 9
rect -19 -5 6 -1
rect 33 -1 37 4
rect 65 8 69 19
rect 84 12 86 16
rect 65 3 69 4
rect 75 8 79 9
rect 11 -5 26 -1
rect 33 -5 49 -1
rect 75 -1 79 4
rect 83 8 87 9
rect 83 -1 87 4
rect 54 -5 68 -1
rect 75 -5 87 -1
rect -19 -9 -15 -5
rect -12 -12 15 -8
rect -12 -15 -7 -12
rect 33 -9 37 -5
rect 75 -9 79 -5
rect 83 -9 87 -5
rect 91 8 95 9
rect 91 0 95 4
rect 99 8 103 19
rect 99 3 103 4
rect 109 8 113 9
rect 109 0 113 4
rect 120 8 124 19
rect 120 3 124 4
rect 130 8 134 9
rect 91 -5 97 0
rect 130 -1 134 4
rect 130 -5 140 -1
rect 91 -9 95 -5
rect 109 -9 113 -5
rect 130 -9 134 -5
rect -19 -20 -12 -16
rect 23 -23 27 -13
rect 45 -20 57 -16
rect 65 -23 69 -13
rect 83 -20 86 -16
rect 99 -23 103 -13
rect 120 -23 124 -13
rect -30 -24 75 -23
rect 92 -24 140 -23
rect -30 -25 140 -24
rect -30 -29 -24 -25
rect -20 -29 35 -25
rect 39 -29 92 -25
rect 96 -29 125 -25
rect 129 -29 140 -25
rect -30 -31 140 -29
rect -30 -42 -26 -31
rect -10 -42 -6 -31
rect 9 -38 21 -34
rect 25 -38 33 -34
rect 41 -42 45 -31
rect 56 -38 79 -34
rect 94 -42 98 -31
rect -36 -55 -27 -51
rect -30 -59 -26 -58
rect -30 -75 -26 -63
rect -20 -59 -16 -46
rect -11 -55 -7 -51
rect -20 -64 -16 -63
rect -10 -59 -6 -58
rect -10 -75 -6 -63
rect 0 -59 4 -46
rect 0 -64 4 -63
rect 18 -58 22 -46
rect 26 -58 30 -46
rect 38 -55 42 -51
rect 76 -52 80 -46
rect 73 -56 80 -52
rect 76 -58 80 -56
rect 102 -42 106 -31
rect 84 -58 88 -46
rect 113 -50 117 -46
rect 95 -55 98 -51
rect 103 -55 106 -51
rect 118 -55 140 -50
rect 113 -58 117 -55
rect 12 -72 21 -68
rect 25 -72 32 -68
rect 41 -75 45 -64
rect 65 -72 79 -68
rect 94 -75 98 -64
rect 102 -75 106 -64
rect -30 -77 127 -75
rect -30 -81 7 -77
rect 11 -81 60 -77
rect 64 -81 98 -77
rect 102 -81 127 -77
rect -30 -83 127 -81
rect 135 -83 138 -75
<< m2contact >>
rect 127 19 135 27
rect -3 11 2 16
rect 6 -5 11 0
rect 79 12 84 17
rect 49 -5 54 0
rect 15 -13 20 -8
rect 97 -5 102 0
rect 109 -5 114 0
rect 118 -5 123 0
rect -12 -20 -7 -15
rect 40 -20 45 -15
rect 57 -20 62 -15
rect 78 -21 83 -16
rect 4 -39 9 -34
rect 33 -39 38 -34
rect 51 -39 56 -34
rect -16 -55 -11 -50
rect 4 -55 9 -50
rect 13 -56 18 -51
rect 42 -55 47 -50
rect 68 -56 73 -51
rect 98 -55 103 -50
rect 113 -55 118 -50
rect 7 -72 12 -67
rect 32 -72 37 -67
rect 60 -72 65 -67
rect 127 -83 135 -75
<< metal2 >>
rect -16 -20 -12 -16
rect -16 -50 -11 -20
rect -3 -34 2 11
rect 15 12 79 16
rect 6 -25 11 -5
rect 15 -8 19 12
rect 33 -20 40 -15
rect 6 -30 18 -25
rect -3 -39 4 -34
rect -3 -40 9 -39
rect 4 -50 9 -40
rect 13 -51 18 -30
rect 33 -34 38 -20
rect 49 -24 53 -5
rect 62 -20 78 -16
rect 66 -24 71 -20
rect 42 -29 53 -24
rect 60 -29 71 -24
rect 97 -25 102 -5
rect 109 -8 114 -5
rect -16 -68 -11 -55
rect 42 -50 47 -29
rect -16 -72 7 -68
rect 52 -68 56 -39
rect 37 -72 56 -68
rect 60 -67 64 -29
rect 78 -31 102 -25
rect 106 -13 114 -8
rect 78 -34 84 -31
rect 68 -39 84 -34
rect 106 -36 111 -13
rect 118 -17 123 -5
rect 68 -51 73 -39
rect 98 -41 111 -36
rect 115 -24 123 -17
rect 98 -50 103 -41
rect 115 -46 120 -24
rect 113 -50 120 -46
rect 118 -51 120 -50
rect 127 -75 135 19
<< labels >>
rlabel metal1 -28 23 -28 23 5 Vdd
rlabel metal1 -28 -27 -28 -27 1 Gnd
rlabel metal1 -28 -1 -28 -1 1 D
rlabel metal1 -28 -53 -28 -53 1 clk
rlabel metal1 137 -3 137 -3 7 Q_bar
rlabel metal1 138 -53 138 -53 7 Q
<< end >>
