magic
tech scmos
timestamp 1480738159
<< nwell >>
rect 154 -101 173 -69
<< pwell >>
rect 32 -132 38 -126
rect 152 -134 171 -102
<< metal1 >>
rect 0 57 5 65
rect 0 39 3 46
rect 0 1 5 9
rect 71 -10 85 -2
rect 0 -28 3 -21
rect 71 -66 85 -58
rect 72 -77 86 -69
rect 154 -77 167 -69
rect 0 -95 3 -88
rect 71 -133 85 -125
rect 153 -133 166 -125
rect 0 -162 3 -155
<< m2contact >>
rect 79 -28 85 -21
rect 80 -95 86 -89
rect 162 -95 167 -88
rect 165 -122 170 -117
<< metal2 >>
rect 72 49 85 54
rect 0 30 3 35
rect 71 -32 75 -13
rect 79 -21 85 49
rect 155 -18 167 -13
rect 0 -37 3 -32
rect 71 -37 84 -32
rect 71 -85 85 -80
rect 80 -89 85 -85
rect 154 -99 158 -80
rect 162 -88 167 -18
rect 234 -85 237 -80
rect 0 -104 3 -99
rect 83 -147 88 -99
rect 154 -104 165 -99
rect 165 -137 170 -122
rect 72 -152 88 -147
rect 0 -171 3 -166
<< m123contact >>
rect 18 58 24 64
rect 2 12 7 17
rect 32 2 38 8
rect 18 -9 24 -3
rect 2 -55 7 -50
rect 97 -55 102 -50
rect 32 -65 38 -59
rect 18 -76 24 -70
rect 2 -122 7 -117
rect 32 -132 38 -126
rect 18 -143 24 -137
rect 97 -122 102 -117
rect 2 -189 7 -184
rect 32 -199 38 -193
<< metal3 >>
rect 2 -50 7 12
rect 2 -117 7 -55
rect 2 -184 7 -122
rect 18 -3 24 58
rect 18 -70 24 -9
rect 18 -137 24 -76
rect 32 -59 38 2
rect 32 -126 38 -65
rect 2 -204 7 -189
rect 32 -193 38 -132
rect 97 -117 102 -55
rect 97 -138 102 -122
use mux21  mux21_0
timestamp 1480737015
transform 1 0 41 0 1 18
box -41 -18 31 47
use mux21  mux21_1
timestamp 1480737015
transform 1 0 41 0 1 -49
box -41 -18 31 47
use mux21  mux21_4
timestamp 1480737015
transform 1 0 124 0 1 -49
box -41 -18 31 47
use mux21  mux21_2
timestamp 1480737015
transform 1 0 41 0 1 -116
box -41 -18 31 47
use mux21  mux21_5
timestamp 1480737015
transform 1 0 124 0 1 -116
box -41 -18 31 47
use mux21  mux21_6
timestamp 1480737015
transform 1 0 206 0 1 -116
box -41 -18 31 47
use mux21  mux21_3
timestamp 1480737015
transform 1 0 41 0 1 -183
box -41 -18 31 47
<< labels >>
rlabel metal2 236 -83 236 -83 7 out
rlabel metal1 1 42 1 42 3 A0
rlabel metal2 1 33 1 33 3 B0
rlabel metal1 1 -25 1 -25 3 A1
rlabel metal2 1 -34 1 -34 3 B1
rlabel metal1 1 -92 1 -92 3 A2
rlabel metal2 1 -101 1 -101 3 B2
rlabel metal1 1 -157 1 -157 3 A3
rlabel metal2 1 -168 1 -168 3 B3
rlabel metal1 2 61 2 61 4 Vdd
rlabel metal1 2 5 2 5 3 Gnd
rlabel metal3 4 -202 4 -202 2 s_input2
rlabel metal3 100 -135 100 -135 1 s_input1
rlabel metal2 167 -135 167 -135 1 s_input0
<< end >>
