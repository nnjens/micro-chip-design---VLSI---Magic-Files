magic
tech scmos
timestamp 1480985955
<< nwell >>
rect -35 1 326 32
<< pwell >>
rect -35 -25 326 1
<< ntransistor >>
rect -24 -10 -22 -5
rect -8 -10 -6 -5
rect 0 -10 2 -5
rect 8 -10 10 -5
rect 24 -10 26 -5
rect 32 -10 34 -5
rect 40 -10 42 -5
rect 48 -10 50 -5
rect 56 -10 58 -5
rect 64 -10 66 -5
rect 72 -10 74 -5
rect 80 -10 82 -5
rect 88 -10 90 -5
rect 104 -10 106 -5
rect 112 -10 114 -5
rect 120 -10 122 -5
rect 128 -10 130 -5
rect 136 -10 138 -5
rect 144 -10 146 -5
rect 152 -10 154 -5
rect 160 -10 162 -5
rect 168 -10 170 -5
rect 176 -10 178 -5
rect 184 -10 186 -5
rect 192 -10 194 -5
rect 200 -10 202 -5
rect 208 -10 210 -5
rect 216 -10 218 -5
rect 224 -10 226 -5
rect 232 -10 234 -5
rect 240 -10 242 -5
rect 248 -10 250 -5
rect 256 -10 258 -5
rect 264 -10 266 -5
rect 272 -10 274 -5
rect 280 -10 282 -5
rect 288 -10 290 -5
rect 296 -10 298 -5
rect 304 -10 306 -5
rect 312 -10 314 -5
<< ptransistor >>
rect -24 7 -22 17
rect -8 7 -6 17
rect 0 7 2 17
rect 8 7 10 17
rect 24 7 26 17
rect 32 7 34 17
rect 40 7 42 17
rect 48 7 50 17
rect 56 7 58 17
rect 64 7 66 17
rect 72 7 74 17
rect 80 7 82 17
rect 88 7 90 17
rect 104 7 106 17
rect 112 7 114 17
rect 120 7 122 17
rect 128 7 130 17
rect 136 7 138 17
rect 144 7 146 17
rect 152 7 154 17
rect 160 7 162 17
rect 168 7 170 17
rect 176 7 178 17
rect 184 7 186 17
rect 192 7 194 17
rect 200 7 202 17
rect 208 7 210 17
rect 216 7 218 17
rect 224 7 226 17
rect 232 7 234 17
rect 240 7 242 17
rect 248 7 250 17
rect 256 7 258 17
rect 264 7 266 17
rect 272 7 274 17
rect 280 7 282 17
rect 288 7 290 17
rect 296 7 298 17
rect 304 7 306 17
rect 312 7 314 17
<< ndiffusion >>
rect -25 -10 -24 -5
rect -22 -10 -21 -5
rect -9 -10 -8 -5
rect -6 -10 0 -5
rect 2 -10 8 -5
rect 10 -10 11 -5
rect 23 -10 24 -5
rect 26 -10 32 -5
rect 34 -10 40 -5
rect 42 -10 48 -5
rect 50 -10 56 -5
rect 58 -10 64 -5
rect 66 -10 72 -5
rect 74 -10 80 -5
rect 82 -10 88 -5
rect 90 -10 91 -5
rect 103 -10 104 -5
rect 106 -10 112 -5
rect 114 -10 120 -5
rect 122 -10 128 -5
rect 130 -10 136 -5
rect 138 -10 144 -5
rect 146 -10 152 -5
rect 154 -10 160 -5
rect 162 -10 168 -5
rect 170 -10 176 -5
rect 178 -10 184 -5
rect 186 -10 192 -5
rect 194 -10 200 -5
rect 202 -10 208 -5
rect 210 -10 216 -5
rect 218 -10 224 -5
rect 226 -10 232 -5
rect 234 -10 240 -5
rect 242 -10 248 -5
rect 250 -10 256 -5
rect 258 -10 264 -5
rect 266 -10 272 -5
rect 274 -10 280 -5
rect 282 -10 288 -5
rect 290 -10 296 -5
rect 298 -10 304 -5
rect 306 -10 312 -5
rect 314 -10 315 -5
<< pdiffusion >>
rect -25 7 -24 17
rect -22 7 -21 17
rect -9 7 -8 17
rect -6 7 -5 17
rect -1 7 0 17
rect 2 7 3 17
rect 7 7 8 17
rect 10 7 11 17
rect 23 7 24 17
rect 26 7 27 17
rect 31 7 32 17
rect 34 7 35 17
rect 39 7 40 17
rect 42 7 43 17
rect 47 7 48 17
rect 50 7 51 17
rect 55 7 56 17
rect 58 7 59 17
rect 63 7 64 17
rect 66 7 67 17
rect 71 7 72 17
rect 74 7 75 17
rect 79 7 80 17
rect 82 7 83 17
rect 87 7 88 17
rect 90 7 91 17
rect 103 7 104 17
rect 106 7 107 17
rect 111 7 112 17
rect 114 7 115 17
rect 119 7 120 17
rect 122 7 123 17
rect 127 7 128 17
rect 130 7 131 17
rect 135 7 136 17
rect 138 7 139 17
rect 143 7 144 17
rect 146 7 147 17
rect 151 7 152 17
rect 154 7 155 17
rect 159 7 160 17
rect 162 7 163 17
rect 167 7 168 17
rect 170 7 171 17
rect 175 7 176 17
rect 178 7 179 17
rect 183 7 184 17
rect 186 7 187 17
rect 191 7 192 17
rect 194 7 195 17
rect 199 7 200 17
rect 202 7 203 17
rect 207 7 208 17
rect 210 7 211 17
rect 215 7 216 17
rect 218 7 219 17
rect 223 7 224 17
rect 226 7 227 17
rect 231 7 232 17
rect 234 7 235 17
rect 239 7 240 17
rect 242 7 243 17
rect 247 7 248 17
rect 250 7 251 17
rect 255 7 256 17
rect 258 7 259 17
rect 263 7 264 17
rect 266 7 267 17
rect 271 7 272 17
rect 274 7 275 17
rect 279 7 280 17
rect 282 7 283 17
rect 287 7 288 17
rect 290 7 291 17
rect 295 7 296 17
rect 298 7 299 17
rect 303 7 304 17
rect 306 7 307 17
rect 311 7 312 17
rect 314 7 315 17
<< ndcontact >>
rect -29 -10 -25 -5
rect -21 -10 -17 -5
rect -13 -10 -9 -5
rect 11 -10 15 -5
rect 19 -10 23 -5
rect 91 -10 95 -5
rect 99 -10 103 -5
rect 315 -10 319 -5
<< pdcontact >>
rect -29 7 -25 17
rect -21 7 -17 17
rect -13 7 -9 17
rect -5 7 -1 17
rect 3 7 7 17
rect 11 7 15 17
rect 19 7 23 17
rect 27 7 31 17
rect 35 7 39 17
rect 43 7 47 17
rect 51 7 55 17
rect 59 7 63 17
rect 67 7 71 17
rect 75 7 79 17
rect 83 7 87 17
rect 91 7 95 17
rect 99 7 103 17
rect 107 7 111 17
rect 115 7 119 17
rect 123 7 127 17
rect 131 7 135 17
rect 139 7 143 17
rect 147 7 151 17
rect 155 7 159 17
rect 163 7 167 17
rect 171 7 175 17
rect 179 7 183 17
rect 187 7 191 17
rect 195 7 199 17
rect 203 7 207 17
rect 211 7 215 17
rect 219 7 223 17
rect 227 7 231 17
rect 235 7 239 17
rect 243 7 247 17
rect 251 7 255 17
rect 259 7 263 17
rect 267 7 271 17
rect 275 7 279 17
rect 283 7 287 17
rect 291 7 295 17
rect 299 7 303 17
rect 307 7 311 17
rect 315 7 319 17
<< polysilicon >>
rect -24 17 -22 20
rect -8 17 -6 20
rect 0 17 2 20
rect 8 17 10 20
rect 24 17 26 20
rect 32 17 34 20
rect 40 17 42 20
rect 48 17 50 20
rect 56 17 58 20
rect 64 17 66 20
rect 72 17 74 20
rect 80 17 82 20
rect 88 17 90 20
rect 104 17 106 20
rect 112 17 114 20
rect 120 17 122 20
rect 128 17 130 20
rect 136 17 138 20
rect 144 17 146 20
rect 152 17 154 20
rect 160 17 162 20
rect 168 17 170 20
rect 176 17 178 20
rect 184 17 186 20
rect 192 17 194 20
rect 200 17 202 20
rect 208 17 210 20
rect 216 17 218 20
rect 224 17 226 20
rect 232 17 234 20
rect 240 17 242 20
rect 248 17 250 20
rect 256 17 258 20
rect 264 17 266 20
rect 272 17 274 20
rect 280 17 282 20
rect 288 17 290 20
rect 296 17 298 20
rect 304 17 306 20
rect 312 17 314 20
rect -24 -5 -22 7
rect -8 3 -6 7
rect 0 3 2 7
rect 8 3 10 7
rect 24 3 26 7
rect 32 3 34 7
rect 40 3 42 7
rect 48 3 50 7
rect 56 3 58 7
rect 64 3 66 7
rect 72 3 74 7
rect 80 3 82 7
rect 88 3 90 7
rect 104 3 106 7
rect 112 3 114 7
rect 120 3 122 7
rect 128 3 130 7
rect 136 3 138 7
rect 144 3 146 7
rect 152 3 154 7
rect 160 3 162 7
rect 168 3 170 7
rect 176 3 178 7
rect 184 3 186 7
rect 192 3 194 7
rect 200 3 202 7
rect 208 3 210 7
rect 216 3 218 7
rect 224 3 226 7
rect 232 3 234 7
rect 240 3 242 7
rect 248 3 250 7
rect 256 3 258 7
rect 264 3 266 7
rect 272 3 274 7
rect 280 3 282 7
rect 288 3 290 7
rect 296 3 298 7
rect 304 3 306 7
rect 312 3 314 7
rect -8 -1 10 3
rect 24 -1 90 3
rect 104 -1 314 3
rect -8 -5 -6 -1
rect 0 -5 2 -1
rect 8 -5 10 -1
rect 24 -5 26 -1
rect 32 -5 34 -1
rect 40 -5 42 -1
rect 48 -5 50 -1
rect 56 -5 58 -1
rect 64 -5 66 -1
rect 72 -5 74 -1
rect 80 -5 82 -1
rect 88 -5 90 -1
rect 104 -5 106 -1
rect 112 -5 114 -1
rect 120 -5 122 -1
rect 128 -5 130 -1
rect 136 -5 138 -1
rect 144 -5 146 -1
rect 152 -5 154 -1
rect 160 -5 162 -1
rect 168 -5 170 -1
rect 176 -5 178 -1
rect 184 -5 186 -1
rect 192 -5 194 -1
rect 200 -5 202 -1
rect 208 -5 210 -1
rect 216 -5 218 -1
rect 224 -5 226 -1
rect 232 -5 234 -1
rect 240 -5 242 -1
rect 248 -5 250 -1
rect 256 -5 258 -1
rect 264 -5 266 -1
rect 272 -5 274 -1
rect 280 -5 282 -1
rect 288 -5 290 -1
rect 296 -5 298 -1
rect 304 -5 306 -1
rect 312 -5 314 -1
rect -24 -13 -22 -10
rect -8 -13 -6 -10
rect 0 -13 2 -10
rect 8 -13 10 -10
rect 24 -13 26 -10
rect 32 -13 34 -10
rect 40 -13 42 -10
rect 48 -13 50 -10
rect 56 -13 58 -10
rect 64 -13 66 -10
rect 72 -13 74 -10
rect 80 -13 82 -10
rect 88 -13 90 -10
rect 104 -13 106 -10
rect 112 -13 114 -10
rect 120 -13 122 -10
rect 128 -13 130 -10
rect 136 -13 138 -10
rect 144 -13 146 -10
rect 152 -13 154 -10
rect 160 -13 162 -10
rect 168 -13 170 -10
rect 176 -13 178 -10
rect 184 -13 186 -10
rect 192 -13 194 -10
rect 200 -13 202 -10
rect 208 -13 210 -10
rect 216 -13 218 -10
rect 224 -13 226 -10
rect 232 -13 234 -10
rect 240 -13 242 -10
rect 248 -13 250 -10
rect 256 -13 258 -10
rect 264 -13 266 -10
rect 272 -13 274 -10
rect 280 -13 282 -10
rect 288 -13 290 -10
rect 296 -13 298 -10
rect 304 -13 306 -10
rect 312 -13 314 -10
<< polycontact >>
rect -28 0 -24 4
rect -12 -1 -8 3
rect 20 -1 24 3
rect 100 -1 104 3
<< metal1 >>
rect -33 23 321 31
rect -29 17 -25 23
rect -13 17 -9 23
rect 3 17 7 23
rect 19 17 23 23
rect 35 17 39 23
rect 51 17 55 23
rect 67 17 71 23
rect 83 17 87 23
rect 99 17 103 23
rect 115 17 119 23
rect 131 17 135 23
rect 147 17 151 23
rect 163 17 167 23
rect 179 17 183 23
rect 195 17 199 23
rect 211 17 215 23
rect 227 17 231 23
rect 243 17 247 23
rect 259 17 263 23
rect 275 17 279 23
rect 291 17 295 23
rect 307 17 311 23
rect -31 0 -28 4
rect -21 3 -17 7
rect -5 3 -1 7
rect 11 3 15 7
rect 27 3 31 7
rect 43 3 47 7
rect 59 3 63 7
rect 75 3 79 7
rect 91 3 95 7
rect 107 3 111 7
rect 123 3 127 7
rect 139 3 143 7
rect 155 3 159 7
rect 171 3 175 7
rect 187 3 191 7
rect 203 3 207 7
rect 219 3 223 7
rect 235 3 239 7
rect 251 3 255 7
rect 267 3 271 7
rect 283 3 287 7
rect 299 3 303 7
rect 315 3 319 7
rect -21 -1 -12 3
rect -5 -1 20 3
rect 27 -1 100 3
rect 107 -1 321 3
rect -21 -5 -17 -1
rect 11 -5 15 -1
rect 91 -5 95 -1
rect 315 -5 319 -1
rect -29 -17 -25 -10
rect -13 -17 -9 -10
rect 19 -17 23 -10
rect 99 -17 103 -10
rect -33 -25 321 -17
<< labels >>
rlabel metal1 -30 26 -30 26 3 Vdd
rlabel metal1 -30 -20 -30 -20 2 Gnd
rlabel metal1 319 1 319 1 1 out
rlabel metal1 -30 2 -30 2 3 in
<< end >>
