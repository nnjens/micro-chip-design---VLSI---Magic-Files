magic
tech scmos
timestamp 1480810385
<< nwell >>
rect -98 405 94 431
rect -98 346 94 375
rect -98 286 94 314
rect -98 227 94 256
rect 69 195 94 197
rect -98 168 94 195
rect -98 135 -65 138
rect -98 109 94 135
rect -98 76 75 77
rect -98 50 94 76
rect -98 -10 94 22
<< pwell >>
rect -98 375 94 405
rect -98 314 94 346
rect -98 256 94 286
rect -98 197 94 227
rect -98 195 69 197
rect -98 143 94 168
rect -98 138 -65 143
rect -98 85 94 109
rect -98 77 75 85
rect -98 22 94 50
rect -98 -34 94 -10
rect -98 -35 75 -34
<< ntransistor >>
rect -83 393 -81 399
rect -43 393 -41 399
rect -23 393 -21 399
rect -3 393 -1 399
rect 15 393 17 399
rect 33 393 35 399
rect 43 393 45 399
rect 60 393 62 399
rect 79 393 81 399
rect -43 334 -41 340
rect -23 334 -21 340
rect -13 334 -11 340
rect 15 334 17 340
rect 33 334 35 340
rect 43 334 45 340
rect 60 334 62 340
rect 79 334 81 340
rect -83 274 -81 280
rect -43 274 -41 280
rect -33 274 -31 280
rect -3 274 -1 280
rect 15 274 17 280
rect 33 274 35 280
rect 43 274 45 280
rect 60 274 62 280
rect 79 274 81 280
rect -43 215 -41 221
rect -33 215 -31 221
rect -13 215 -11 221
rect 15 215 17 221
rect 33 215 35 221
rect 43 215 45 221
rect 60 215 62 221
rect 79 215 81 221
rect -83 156 -81 162
rect -53 156 -51 162
rect -53 97 -51 103
rect -79 38 -77 44
rect -71 38 -69 44
rect -53 38 -51 44
rect -77 -22 -75 -16
rect -53 -22 -51 -16
rect -23 156 -21 162
rect -3 156 -1 162
rect 15 156 17 162
rect 33 156 35 162
rect 43 156 45 162
rect 60 156 62 162
rect 79 156 81 162
rect -23 97 -21 103
rect -13 97 -11 103
rect -33 38 -31 44
rect -33 -22 -31 -16
rect 14 97 16 103
rect 33 97 35 103
rect 43 97 45 103
rect 60 97 62 103
rect 79 97 81 103
rect -3 38 -1 44
rect 15 38 17 44
rect 33 38 35 44
rect 43 38 45 44
rect 60 38 62 44
rect 79 38 81 44
rect -13 -22 -11 -16
rect 14 -22 16 -16
rect 33 -22 35 -16
rect 43 -22 45 -16
rect 60 -22 62 -16
rect 79 -22 81 -16
<< ptransistor >>
rect -83 411 -81 419
rect -43 411 -41 419
rect -23 411 -21 419
rect -3 411 -1 419
rect 15 411 17 419
rect 33 411 35 419
rect 43 411 45 419
rect 60 411 62 419
rect 79 411 81 419
rect -43 352 -41 360
rect -23 352 -21 360
rect -13 352 -11 360
rect 15 352 17 360
rect 33 352 35 360
rect 43 352 45 360
rect 60 352 62 360
rect 79 352 81 360
rect -83 292 -81 300
rect -43 292 -41 300
rect -33 292 -31 300
rect -3 292 -1 300
rect 15 292 17 300
rect 33 292 35 300
rect 43 292 45 300
rect 60 292 62 300
rect 79 292 81 300
rect -43 233 -41 241
rect -33 233 -31 241
rect -13 233 -11 241
rect 15 233 17 241
rect 33 233 35 241
rect 43 233 45 241
rect 60 233 62 241
rect 79 233 81 241
rect -83 174 -81 182
rect -53 174 -51 182
rect -53 115 -51 123
rect -79 56 -77 64
rect -71 56 -69 64
rect -53 56 -51 64
rect -77 -4 -75 4
rect -53 -4 -51 4
rect -23 174 -21 182
rect -3 174 -1 182
rect 15 174 17 182
rect 33 174 35 182
rect 43 174 45 182
rect 60 174 62 182
rect 79 174 81 182
rect -23 115 -21 123
rect -13 115 -11 123
rect -33 56 -31 64
rect -33 -4 -31 4
rect 14 115 16 123
rect 33 115 35 123
rect 43 115 45 123
rect 60 115 62 123
rect 79 115 81 123
rect -3 56 -1 64
rect 15 56 17 64
rect 33 56 35 64
rect 43 56 45 64
rect 60 56 62 64
rect 79 56 81 64
rect -13 -4 -11 4
rect 14 -4 16 4
rect 33 -4 35 4
rect 43 -4 45 4
rect 60 -4 62 4
rect 79 -4 81 4
<< ndiffusion >>
rect -85 393 -83 399
rect -81 393 -78 399
rect -45 393 -43 399
rect -41 393 -39 399
rect -25 393 -23 399
rect -21 393 -19 399
rect -5 393 -3 399
rect -1 393 1 399
rect 13 393 15 399
rect 17 393 20 399
rect 32 393 33 399
rect 35 393 43 399
rect 45 393 46 399
rect 58 393 60 399
rect 62 393 65 399
rect 77 393 79 399
rect 81 393 84 399
rect -45 334 -43 340
rect -41 334 -39 340
rect -25 334 -23 340
rect -21 334 -13 340
rect -11 334 -10 340
rect 13 334 15 340
rect 17 334 20 340
rect 32 334 33 340
rect 35 334 43 340
rect 45 334 46 340
rect 58 334 60 340
rect 62 334 65 340
rect 77 334 79 340
rect 81 334 84 340
rect -85 274 -83 280
rect -81 274 -78 280
rect -45 274 -43 280
rect -41 274 -33 280
rect -31 274 -30 280
rect -5 274 -3 280
rect -1 274 0 280
rect 13 274 15 280
rect 17 274 20 280
rect 32 274 33 280
rect 35 274 43 280
rect 45 274 46 280
rect 58 274 60 280
rect 62 274 65 280
rect 77 274 79 280
rect 81 274 84 280
rect -45 215 -43 221
rect -41 215 -33 221
rect -31 215 -30 221
rect -15 215 -13 221
rect -11 215 -10 221
rect 13 215 15 221
rect 17 215 20 221
rect 32 215 33 221
rect 35 215 43 221
rect 45 215 46 221
rect 58 215 60 221
rect 62 215 65 221
rect 77 215 79 221
rect 81 215 84 221
rect -85 156 -83 162
rect -81 156 -78 162
rect -55 156 -53 162
rect -51 156 -49 162
rect -55 97 -53 103
rect -51 97 -49 103
rect -80 38 -79 44
rect -77 38 -76 44
rect -72 38 -71 44
rect -69 38 -68 44
rect -55 38 -53 44
rect -51 38 -49 44
rect -79 -22 -77 -16
rect -75 -22 -72 -16
rect -55 -22 -53 -16
rect -51 -22 -49 -16
rect -26 156 -23 162
rect -21 156 -20 162
rect -5 156 -3 162
rect -1 156 1 162
rect 13 156 15 162
rect 17 156 20 162
rect 32 156 33 162
rect 35 156 43 162
rect 45 156 46 162
rect 58 156 60 162
rect 62 156 65 162
rect 77 156 79 162
rect 81 156 84 162
rect -25 97 -23 103
rect -21 97 -13 103
rect -11 97 -9 103
rect -35 38 -33 44
rect -31 38 -29 44
rect -35 -22 -33 -16
rect -31 -22 -29 -16
rect 12 97 14 103
rect 16 97 19 103
rect 32 97 33 103
rect 35 97 43 103
rect 45 97 46 103
rect 58 97 60 103
rect 62 97 65 103
rect 77 97 79 103
rect 81 97 84 103
rect -5 38 -3 44
rect -1 38 1 44
rect 13 38 15 44
rect 17 38 20 44
rect 32 38 33 44
rect 35 38 43 44
rect 45 38 46 44
rect 58 38 60 44
rect 62 38 65 44
rect 77 38 79 44
rect 81 38 84 44
rect -15 -22 -13 -16
rect -11 -22 -9 -16
rect 12 -22 14 -16
rect 16 -22 19 -16
rect 32 -22 33 -16
rect 35 -22 43 -16
rect 45 -22 46 -16
rect 58 -22 60 -16
rect 62 -22 65 -16
rect 77 -22 79 -16
rect 81 -22 84 -16
<< pdiffusion >>
rect -85 411 -83 419
rect -81 411 -78 419
rect -45 411 -43 419
rect -41 411 -39 419
rect -25 411 -23 419
rect -21 411 -18 419
rect -5 411 -3 419
rect -1 411 1 419
rect 13 411 15 419
rect 17 411 20 419
rect 32 411 33 419
rect 35 411 38 419
rect 42 411 43 419
rect 45 411 46 419
rect 58 411 60 419
rect 62 411 65 419
rect 77 411 79 419
rect 81 411 84 419
rect -45 352 -43 360
rect -41 352 -39 360
rect -25 352 -23 360
rect -21 352 -19 360
rect -15 352 -13 360
rect -11 352 -10 360
rect 13 352 15 360
rect 17 352 20 360
rect 32 352 33 360
rect 35 352 38 360
rect 42 352 43 360
rect 45 352 46 360
rect 58 352 60 360
rect 62 352 65 360
rect 77 352 79 360
rect 81 352 84 360
rect -85 292 -83 300
rect -81 292 -78 300
rect -45 292 -43 300
rect -41 292 -39 300
rect -35 292 -33 300
rect -31 292 -29 300
rect -5 292 -3 300
rect -1 292 1 300
rect 13 292 15 300
rect 17 292 20 300
rect 32 292 33 300
rect 35 292 38 300
rect 42 292 43 300
rect 45 292 46 300
rect 58 292 60 300
rect 62 292 65 300
rect 77 292 79 300
rect 81 292 84 300
rect -45 233 -43 241
rect -41 233 -39 241
rect -35 233 -33 241
rect -31 233 -29 241
rect -15 233 -13 241
rect -11 233 -9 241
rect 13 233 15 241
rect 17 233 20 241
rect 32 233 33 241
rect 35 233 38 241
rect 42 233 43 241
rect 45 233 46 241
rect 58 233 60 241
rect 62 233 65 241
rect 77 233 79 241
rect 81 233 84 241
rect -85 174 -83 182
rect -81 174 -78 182
rect -55 174 -53 182
rect -51 174 -49 182
rect -55 115 -53 123
rect -51 115 -49 123
rect -80 56 -79 64
rect -77 56 -76 64
rect -72 56 -71 64
rect -69 56 -68 64
rect -55 56 -53 64
rect -51 56 -49 64
rect -79 -4 -77 4
rect -75 -4 -72 4
rect -55 -4 -53 4
rect -51 -4 -49 4
rect -26 174 -23 182
rect -21 174 -20 182
rect -5 174 -3 182
rect -1 174 1 182
rect 13 174 15 182
rect 17 174 20 182
rect 32 174 33 182
rect 35 174 38 182
rect 42 174 43 182
rect 45 174 46 182
rect 58 174 60 182
rect 62 174 65 182
rect 77 174 79 182
rect 81 174 84 182
rect -25 115 -23 123
rect -21 115 -19 123
rect -15 115 -13 123
rect -11 115 -9 123
rect -35 56 -33 64
rect -31 56 -29 64
rect -35 -4 -33 4
rect -31 -4 -29 4
rect 12 115 14 123
rect 16 115 19 123
rect 32 115 33 123
rect 35 115 38 123
rect 42 115 43 123
rect 45 115 46 123
rect 58 115 60 123
rect 62 115 65 123
rect 77 115 79 123
rect 81 115 84 123
rect -5 56 -3 64
rect -1 56 1 64
rect 13 56 15 64
rect 17 56 20 64
rect 32 56 33 64
rect 35 56 38 64
rect 42 56 43 64
rect 45 56 46 64
rect 58 56 60 64
rect 62 56 65 64
rect 77 56 79 64
rect 81 56 84 64
rect -15 -4 -13 4
rect -11 -4 -9 4
rect 12 -4 14 4
rect 16 -4 19 4
rect 32 -4 33 4
rect 35 -4 38 4
rect 42 -4 43 4
rect 45 -4 46 4
rect 58 -4 60 4
rect 62 -4 65 4
rect 77 -4 79 4
rect 81 -4 84 4
<< ndcontact >>
rect -89 393 -85 399
rect -78 393 -74 399
rect -49 393 -45 399
rect -39 393 -35 399
rect -29 393 -25 399
rect -19 393 -15 399
rect -9 393 -5 399
rect 1 393 5 399
rect 9 393 13 399
rect 20 393 24 399
rect 28 393 32 399
rect 46 393 50 399
rect 54 393 58 399
rect 65 393 69 399
rect 73 393 77 399
rect 84 393 88 399
rect -49 334 -45 340
rect -39 334 -35 340
rect -29 334 -25 340
rect -10 334 -6 340
rect 9 334 13 340
rect 20 334 24 340
rect 28 334 32 340
rect 46 334 50 340
rect 54 334 58 340
rect 65 334 69 340
rect 73 334 77 340
rect 84 334 88 340
rect -89 274 -85 280
rect -78 274 -74 280
rect -49 274 -45 280
rect -30 274 -26 280
rect -9 274 -5 280
rect 0 274 4 280
rect 9 274 13 280
rect 20 274 24 280
rect 28 274 32 280
rect 46 274 50 280
rect 54 274 58 280
rect 65 274 69 280
rect 73 274 77 280
rect 84 274 88 280
rect -49 215 -45 221
rect -30 215 -26 221
rect -19 215 -15 221
rect -10 215 -6 221
rect 9 215 13 221
rect 20 215 24 221
rect 28 215 32 221
rect 46 215 50 221
rect 54 215 58 221
rect 65 215 69 221
rect 73 215 77 221
rect 84 215 88 221
rect -89 156 -85 162
rect -78 156 -74 162
rect -59 156 -55 162
rect -49 156 -45 162
rect -59 97 -55 103
rect -49 97 -45 103
rect -84 38 -80 44
rect -76 38 -72 44
rect -68 38 -64 44
rect -59 38 -55 44
rect -49 38 -45 44
rect -83 -22 -79 -16
rect -72 -22 -68 -16
rect -59 -22 -55 -16
rect -49 -22 -45 -16
rect -30 156 -26 162
rect -20 156 -16 162
rect -9 156 -5 162
rect 1 156 5 162
rect 9 156 13 162
rect 20 156 24 162
rect 28 156 32 162
rect 46 156 50 162
rect 54 156 58 162
rect 65 156 69 162
rect 73 156 77 162
rect 84 156 88 162
rect -29 97 -25 103
rect -9 97 -5 103
rect -39 38 -35 44
rect -29 38 -25 44
rect -39 -22 -35 -16
rect -29 -22 -25 -16
rect 8 97 12 103
rect 19 97 23 103
rect 28 97 32 103
rect 46 97 50 103
rect 54 97 58 103
rect 65 97 69 103
rect 73 97 77 103
rect 84 97 88 103
rect -9 38 -5 44
rect 1 38 5 44
rect 9 38 13 44
rect 20 38 24 44
rect 28 38 32 44
rect 46 38 50 44
rect 54 38 58 44
rect 65 38 69 44
rect 73 38 77 44
rect 84 38 88 44
rect -19 -22 -15 -16
rect -9 -22 -5 -16
rect 8 -22 12 -16
rect 19 -22 23 -16
rect 28 -22 32 -16
rect 46 -22 50 -16
rect 54 -22 58 -16
rect 65 -22 69 -16
rect 73 -22 77 -16
rect 84 -22 88 -16
<< pdcontact >>
rect -89 411 -85 419
rect -78 411 -74 419
rect -49 411 -45 419
rect -39 411 -35 419
rect -29 411 -25 419
rect -18 411 -14 419
rect -9 411 -5 419
rect 1 411 5 419
rect 9 411 13 419
rect 20 411 24 419
rect 28 411 32 419
rect 38 411 42 419
rect 46 411 50 419
rect 54 411 58 419
rect 65 411 69 419
rect 73 411 77 419
rect 84 411 88 419
rect -49 352 -45 360
rect -39 352 -35 360
rect -29 352 -25 360
rect -19 352 -15 360
rect -10 352 -6 360
rect 9 352 13 360
rect 20 352 24 360
rect 28 352 32 360
rect 38 352 42 360
rect 46 352 50 360
rect 54 352 58 360
rect 65 352 69 360
rect 73 352 77 360
rect 84 352 88 360
rect -89 292 -85 300
rect -78 292 -74 300
rect -49 292 -45 300
rect -39 292 -35 300
rect -29 292 -25 300
rect -9 292 -5 300
rect 1 292 5 300
rect 9 292 13 300
rect 20 292 24 300
rect 28 292 32 300
rect 38 292 42 300
rect 46 292 50 300
rect 54 292 58 300
rect 65 292 69 300
rect 73 292 77 300
rect 84 292 88 300
rect -49 233 -45 241
rect -39 233 -35 241
rect -29 233 -25 241
rect -19 233 -15 241
rect -9 233 -5 241
rect 9 233 13 241
rect 20 233 24 241
rect 28 233 32 241
rect 38 233 42 241
rect 46 233 50 241
rect 54 233 58 241
rect 65 233 69 241
rect 73 233 77 241
rect 84 233 88 241
rect -89 174 -85 182
rect -78 174 -74 182
rect -59 174 -55 182
rect -49 174 -45 182
rect -59 115 -55 123
rect -49 115 -45 123
rect -84 56 -80 64
rect -76 56 -72 64
rect -68 56 -64 64
rect -59 56 -55 64
rect -49 56 -45 64
rect -83 -4 -79 4
rect -72 -4 -68 4
rect -59 -4 -55 4
rect -49 -4 -45 4
rect -30 174 -26 182
rect -20 174 -16 182
rect -9 174 -5 182
rect 1 174 5 182
rect 9 174 13 182
rect 20 174 24 182
rect 28 174 32 182
rect 38 174 42 182
rect 46 174 50 182
rect 54 174 58 182
rect 65 174 69 182
rect 73 174 77 182
rect 84 174 88 182
rect -29 115 -25 123
rect -19 115 -15 123
rect -9 115 -5 123
rect -39 56 -35 64
rect -29 56 -25 64
rect -39 -4 -35 4
rect -29 -4 -25 4
rect 8 115 12 123
rect 19 115 23 123
rect 28 115 32 123
rect 38 115 42 123
rect 46 115 50 123
rect 54 115 58 123
rect 65 115 69 123
rect 73 115 77 123
rect 84 115 88 123
rect -9 56 -5 64
rect 1 56 5 64
rect 9 56 13 64
rect 20 56 24 64
rect 28 56 32 64
rect 38 56 42 64
rect 46 56 50 64
rect 54 56 58 64
rect 65 56 69 64
rect 73 56 77 64
rect 84 56 88 64
rect -19 -4 -15 4
rect -9 -4 -5 4
rect 8 -4 12 4
rect 19 -4 23 4
rect 28 -4 32 4
rect 38 -4 42 4
rect 46 -4 50 4
rect 54 -4 58 4
rect 65 -4 69 4
rect 73 -4 77 4
rect 84 -4 88 4
<< psubstratepcontact >>
rect -83 383 -79 387
rect -49 383 -45 387
rect 15 383 19 387
rect 59 383 63 387
rect -49 324 -45 328
rect -83 264 -79 268
rect -49 264 -45 268
rect 15 324 19 328
rect 59 324 63 328
rect 15 264 19 268
rect 59 264 63 268
rect -49 205 -45 209
rect -83 146 -79 150
rect -49 146 -45 150
rect -49 87 -45 91
rect -49 28 -45 32
rect -49 -32 -45 -28
rect 15 205 19 209
rect 59 205 63 209
rect 15 146 19 150
rect 60 146 64 150
rect 13 87 17 91
rect 59 87 63 91
rect 15 28 19 32
rect 60 28 64 32
rect 13 -32 17 -28
rect 59 -32 63 -28
<< nsubstratencontact >>
rect -84 424 -80 428
rect -49 424 -45 428
rect 14 424 18 428
rect 62 424 66 428
rect -49 365 -45 369
rect 14 365 18 369
rect 62 365 66 369
rect -84 305 -80 309
rect -49 305 -45 309
rect -49 246 -45 250
rect 14 305 18 309
rect 62 305 66 309
rect 14 246 18 250
rect 62 246 66 250
rect -84 187 -80 191
rect -49 187 -45 191
rect -49 128 -45 132
rect -49 69 -45 73
rect -49 9 -45 13
rect 15 187 19 191
rect 61 187 65 191
rect 14 128 18 132
rect 61 128 65 132
rect 15 69 19 73
rect 61 69 65 73
rect 14 9 18 13
rect 61 9 65 13
<< polysilicon >>
rect -83 419 -81 422
rect -53 419 -51 431
rect -43 419 -41 431
rect -33 419 -31 431
rect -23 419 -21 431
rect -13 419 -11 431
rect -3 419 -1 431
rect 15 419 17 422
rect 33 419 35 422
rect 43 419 45 431
rect 60 419 62 422
rect 79 419 81 422
rect -83 408 -81 411
rect -83 399 -81 404
rect -53 399 -51 411
rect -43 399 -41 411
rect -33 399 -31 411
rect -23 399 -21 411
rect -13 399 -11 411
rect -3 399 -1 411
rect 15 408 17 411
rect 33 408 35 411
rect 15 399 17 404
rect 33 399 35 404
rect 43 399 45 411
rect 60 408 62 411
rect 79 408 81 411
rect 60 399 62 404
rect 79 399 81 404
rect -83 390 -81 393
rect -53 378 -51 393
rect -53 360 -51 374
rect -43 360 -41 393
rect -33 360 -31 393
rect -23 360 -21 393
rect -13 360 -11 393
rect -3 360 -1 393
rect 15 390 17 393
rect 33 390 35 393
rect 15 360 17 363
rect 33 360 35 363
rect 43 360 45 393
rect 60 390 62 393
rect 79 390 81 393
rect 60 360 62 363
rect 79 360 81 363
rect -53 340 -51 352
rect -43 340 -41 352
rect -33 340 -31 352
rect -23 340 -21 352
rect -13 340 -11 352
rect -3 340 -1 352
rect 15 349 17 352
rect 33 349 35 352
rect 15 340 17 345
rect 33 340 35 345
rect 43 340 45 352
rect 60 349 62 352
rect 79 349 81 352
rect 60 340 62 345
rect 79 340 81 345
rect -83 300 -81 303
rect -53 300 -51 334
rect -43 319 -41 334
rect -43 300 -41 315
rect -33 300 -31 334
rect -23 300 -21 334
rect -83 289 -81 292
rect -83 280 -81 285
rect -53 280 -51 292
rect -43 280 -41 292
rect -33 280 -31 292
rect -23 280 -21 292
rect -83 271 -81 274
rect -53 241 -51 274
rect -43 241 -41 274
rect -33 259 -31 274
rect -33 241 -31 255
rect -23 241 -21 274
rect -13 300 -11 334
rect -3 300 -1 334
rect 15 331 17 334
rect 33 331 35 334
rect 15 300 17 303
rect 33 300 35 303
rect 43 300 45 334
rect 60 331 62 334
rect 79 331 81 334
rect 60 300 62 303
rect 79 300 81 303
rect -13 280 -11 292
rect -3 280 -1 292
rect 15 289 17 292
rect 33 289 35 292
rect 15 280 17 285
rect 33 280 35 285
rect 43 280 45 292
rect 60 289 62 292
rect 79 289 81 292
rect 60 280 62 285
rect 79 280 81 285
rect -13 241 -11 274
rect -3 241 -1 274
rect 15 271 17 274
rect 33 271 35 274
rect 15 241 17 244
rect 33 241 35 244
rect 43 241 45 274
rect 60 271 62 274
rect 79 271 81 274
rect 60 241 62 244
rect 79 241 81 244
rect -53 221 -51 233
rect -43 221 -41 233
rect -33 221 -31 233
rect -23 221 -21 233
rect -13 221 -11 233
rect -3 221 -1 233
rect 15 230 17 233
rect 33 230 35 233
rect 15 221 17 226
rect 33 221 35 226
rect 43 221 45 233
rect 60 230 62 233
rect 79 230 81 233
rect 60 221 62 226
rect 79 221 81 226
rect -83 182 -81 185
rect -53 182 -51 215
rect -83 171 -81 174
rect -83 162 -81 167
rect -53 162 -51 174
rect -83 153 -81 156
rect -53 123 -51 156
rect -53 103 -51 115
rect -88 70 -69 72
rect -79 64 -77 67
rect -71 64 -69 70
rect -53 64 -51 97
rect -79 44 -77 56
rect -71 44 -69 56
rect -53 44 -51 56
rect -79 34 -77 38
rect -71 34 -69 38
rect -77 4 -75 7
rect -53 4 -51 38
rect -77 -7 -75 -4
rect -77 -16 -75 -11
rect -53 -16 -51 -4
rect -77 -25 -75 -22
rect -53 -34 -51 -22
rect -43 -34 -41 215
rect -33 182 -31 215
rect -23 200 -21 215
rect -23 182 -21 196
rect -13 182 -11 215
rect -3 182 -1 215
rect 15 212 17 215
rect 33 212 35 215
rect 15 182 17 185
rect 33 182 35 185
rect 43 182 45 215
rect 60 212 62 215
rect 79 212 81 215
rect 60 182 62 185
rect 79 182 81 185
rect -33 162 -31 174
rect -23 162 -21 174
rect -13 162 -11 174
rect -3 162 -1 174
rect 15 171 17 174
rect 33 171 35 174
rect 15 162 17 167
rect 33 162 35 167
rect 43 162 45 174
rect 60 171 62 174
rect 79 171 81 174
rect 60 162 62 167
rect 79 162 81 167
rect -33 123 -31 156
rect -23 123 -21 156
rect -13 141 -11 156
rect -13 123 -11 137
rect -33 103 -31 115
rect -23 103 -21 115
rect -13 103 -11 115
rect -33 64 -31 97
rect -33 44 -31 56
rect -33 4 -31 38
rect -33 -16 -31 -4
rect -33 -34 -31 -22
rect -23 -34 -21 97
rect -13 64 -11 97
rect -3 82 -1 156
rect 15 153 17 156
rect 33 153 35 156
rect 14 123 16 126
rect 33 123 35 126
rect 43 123 45 156
rect 60 153 62 156
rect 79 153 81 156
rect 60 123 62 126
rect 79 123 81 126
rect 14 112 16 115
rect 33 112 35 115
rect 14 103 16 108
rect 33 103 35 108
rect 43 103 45 115
rect 60 112 62 115
rect 79 112 81 115
rect 60 103 62 108
rect 79 103 81 108
rect 14 94 16 97
rect 33 94 35 97
rect -3 64 -1 78
rect 15 64 17 67
rect 33 64 35 67
rect 43 64 45 97
rect 60 94 62 97
rect 79 94 81 97
rect 60 64 62 67
rect 79 64 81 67
rect -13 44 -11 56
rect -3 44 -1 56
rect 15 53 17 56
rect 33 53 35 56
rect 15 44 17 49
rect 33 44 35 49
rect 43 44 45 56
rect 60 53 62 56
rect 79 53 81 56
rect 60 44 62 49
rect 79 44 81 49
rect -13 4 -11 38
rect -13 -16 -11 -4
rect -13 -34 -11 -22
rect -3 -34 -1 38
rect 15 35 17 38
rect 33 35 35 38
rect 43 23 45 38
rect 60 35 62 38
rect 79 35 81 38
rect 14 4 16 7
rect 33 4 35 7
rect 43 4 45 19
rect 60 4 62 7
rect 79 4 81 7
rect 14 -7 16 -4
rect 33 -7 35 -4
rect 14 -16 16 -11
rect 33 -16 35 -11
rect 43 -16 45 -4
rect 60 -7 62 -4
rect 79 -7 81 -4
rect 60 -16 62 -11
rect 79 -16 81 -11
rect 14 -25 16 -22
rect 33 -25 35 -22
rect 43 -34 45 -22
rect 60 -25 62 -22
rect 79 -25 81 -22
<< polycontact >>
rect -85 404 -81 408
rect 13 404 17 408
rect 31 404 35 408
rect 58 404 62 408
rect 77 404 81 408
rect -55 374 -51 378
rect 13 345 17 349
rect 31 345 35 349
rect 58 345 62 349
rect 77 345 81 349
rect -45 315 -41 319
rect -85 285 -81 289
rect -35 255 -31 259
rect 13 285 17 289
rect 31 285 35 289
rect 58 285 62 289
rect 77 285 81 289
rect 13 226 17 230
rect 31 226 35 230
rect 58 226 62 230
rect 77 226 81 230
rect -85 167 -81 171
rect -92 70 -88 74
rect -83 47 -79 51
rect -79 -11 -75 -7
rect -25 196 -21 200
rect 13 167 17 171
rect 31 167 35 171
rect 58 167 62 171
rect 77 167 81 171
rect -15 137 -11 141
rect 12 108 16 112
rect 31 108 35 112
rect 58 108 62 112
rect 77 108 81 112
rect -5 78 -1 82
rect 13 49 17 53
rect 31 49 35 53
rect 58 49 62 53
rect 77 49 81 53
rect 41 19 45 23
rect 12 -11 16 -7
rect 31 -11 35 -7
rect 58 -11 62 -7
rect 77 -11 81 -7
<< polypplus >>
rect -53 411 -51 419
rect -33 411 -31 419
rect -13 411 -11 419
rect -53 352 -51 360
rect -33 352 -31 360
rect -3 352 -1 360
rect -53 292 -51 300
rect -23 292 -21 300
rect -13 292 -11 300
rect -53 233 -51 241
rect -23 233 -21 241
rect -3 233 -1 241
rect -33 174 -31 182
rect -13 174 -11 182
rect -33 115 -31 123
rect -13 56 -11 64
<< polynplus >>
rect -53 393 -51 399
rect -33 393 -31 399
rect -13 393 -11 399
rect -53 334 -51 340
rect -33 334 -31 340
rect -3 334 -1 340
rect -53 274 -51 280
rect -23 274 -21 280
rect -13 274 -11 280
rect -53 215 -51 221
rect -23 215 -21 221
rect -3 215 -1 221
rect -33 156 -31 162
rect -13 156 -11 162
rect -33 97 -31 103
rect -13 38 -11 44
<< metal1 >>
rect -89 428 21 430
rect -89 424 -84 428
rect -80 424 -49 428
rect -45 424 14 428
rect 18 424 21 428
rect -89 422 21 424
rect 29 428 88 430
rect 29 424 62 428
rect 66 424 88 428
rect 29 422 88 424
rect -89 419 -85 422
rect -59 419 -55 422
rect -18 419 -14 422
rect 9 419 13 422
rect 28 419 32 422
rect 46 419 50 422
rect -59 411 -49 419
rect -35 411 -29 419
rect -14 411 -9 419
rect 54 419 58 422
rect 73 419 77 422
rect -98 404 -85 408
rect -97 319 -93 404
rect -78 399 -74 411
rect -29 408 -25 411
rect 1 408 5 411
rect 20 408 24 411
rect 38 408 42 411
rect 65 408 69 411
rect 84 408 94 411
rect -29 404 13 408
rect 20 404 31 408
rect 38 404 58 408
rect 65 404 77 408
rect 1 399 5 404
rect 20 399 24 404
rect 46 399 50 404
rect 84 399 88 408
rect -59 393 -49 399
rect -35 393 -29 399
rect -15 393 -9 399
rect -89 389 -85 393
rect -59 389 -55 393
rect 9 389 13 393
rect 28 389 32 393
rect 54 389 58 393
rect 73 389 77 393
rect -89 387 43 389
rect -89 383 -83 387
rect -79 383 -49 387
rect -45 383 15 387
rect 19 383 43 387
rect -89 381 43 383
rect 52 387 87 389
rect 52 383 59 387
rect 63 383 87 387
rect 52 381 87 383
rect -69 374 -55 378
rect -65 369 21 371
rect -65 365 -49 369
rect -45 365 14 369
rect 18 365 21 369
rect -65 363 21 365
rect 29 369 88 371
rect 29 365 62 369
rect 66 365 88 369
rect 29 363 88 365
rect -59 360 -55 363
rect -19 360 -15 363
rect 9 360 13 363
rect 28 360 32 363
rect 46 360 50 363
rect -59 352 -49 360
rect -35 352 -29 360
rect 54 360 58 363
rect 73 360 77 363
rect -29 349 -25 352
rect -10 349 -6 352
rect 20 349 24 352
rect 38 349 42 352
rect 65 349 69 352
rect 84 349 94 352
rect -29 345 13 349
rect 20 345 31 349
rect 38 345 58 349
rect 65 345 77 349
rect -10 340 -6 345
rect 20 340 24 345
rect 46 340 50 345
rect 84 340 88 349
rect -59 334 -49 340
rect -35 334 -29 340
rect -59 330 -55 334
rect 9 330 13 334
rect 28 330 32 334
rect 54 330 58 334
rect 73 330 77 334
rect -62 328 43 330
rect -62 324 -49 328
rect -45 324 15 328
rect 19 324 43 328
rect -62 322 43 324
rect 52 328 87 330
rect 52 324 59 328
rect 63 324 87 328
rect 52 322 87 324
rect -97 315 -45 319
rect -89 309 21 311
rect -89 305 -84 309
rect -80 305 -49 309
rect -45 305 14 309
rect 18 305 21 309
rect -89 303 21 305
rect 29 309 88 311
rect 29 305 62 309
rect 66 305 88 309
rect 29 303 88 305
rect -89 300 -85 303
rect -59 300 -55 303
rect -29 300 -25 303
rect 9 300 13 303
rect 28 300 32 303
rect 46 300 50 303
rect -59 292 -49 300
rect -25 292 -9 300
rect 54 300 58 303
rect 73 300 77 303
rect -98 285 -85 289
rect -97 200 -93 285
rect -78 280 -74 292
rect -39 289 -35 292
rect 1 289 5 292
rect 20 289 24 292
rect 38 289 42 292
rect 65 289 69 292
rect 84 289 94 292
rect -39 285 13 289
rect 20 285 31 289
rect 38 285 58 289
rect 65 285 77 289
rect 0 280 4 285
rect 20 280 24 285
rect 46 280 50 285
rect 84 280 88 289
rect -59 274 -49 280
rect -26 274 -9 280
rect -89 270 -85 274
rect -59 270 -55 274
rect 9 270 13 274
rect 28 270 32 274
rect 54 270 58 274
rect 73 270 77 274
rect -89 268 43 270
rect -89 264 -83 268
rect -79 264 -49 268
rect -45 264 15 268
rect 19 264 43 268
rect -89 262 43 264
rect 52 268 87 270
rect 52 264 59 268
rect 63 264 87 268
rect 52 262 87 264
rect -69 255 -35 259
rect -65 250 21 252
rect -65 246 -49 250
rect -45 246 14 250
rect 18 246 21 250
rect -65 244 21 246
rect 29 250 88 252
rect 29 246 62 250
rect 66 246 88 250
rect 29 244 88 246
rect -59 241 -55 244
rect -29 241 -25 244
rect 9 241 13 244
rect 28 241 32 244
rect 46 241 50 244
rect -59 233 -49 241
rect -25 233 -19 241
rect 54 241 58 244
rect 73 241 77 244
rect -39 230 -35 233
rect -9 230 -5 233
rect 20 230 24 233
rect 38 230 42 233
rect 65 230 69 233
rect 84 230 94 233
rect -39 226 13 230
rect 20 226 31 230
rect 38 226 58 230
rect 65 226 77 230
rect -10 221 -6 226
rect 20 221 24 226
rect 46 221 50 226
rect 84 221 88 230
rect -59 215 -49 221
rect -26 215 -19 221
rect -59 211 -55 215
rect 9 211 13 215
rect 28 211 32 215
rect 54 211 58 215
rect 73 211 77 215
rect -62 209 43 211
rect -62 205 -49 209
rect -45 205 15 209
rect 19 205 43 209
rect -62 203 43 205
rect 52 209 87 211
rect 52 205 59 209
rect 63 205 87 209
rect 52 203 87 205
rect -97 196 -25 200
rect -89 191 21 193
rect -89 187 -84 191
rect -80 187 -49 191
rect -45 187 15 191
rect 19 187 21 191
rect -89 185 21 187
rect 29 191 88 193
rect 29 187 61 191
rect 65 187 88 191
rect 29 185 88 187
rect -89 182 -85 185
rect -59 182 -55 185
rect -20 182 -16 185
rect 9 182 13 185
rect 28 182 32 185
rect 46 182 50 185
rect -45 174 -30 182
rect -16 174 -9 182
rect 54 182 58 185
rect 73 182 77 185
rect -98 167 -85 171
rect -97 82 -93 167
rect -78 162 -74 174
rect -30 171 -26 174
rect 1 171 5 174
rect 20 171 24 174
rect 38 171 42 174
rect 65 171 69 174
rect 84 171 94 174
rect -30 167 13 171
rect 20 167 31 171
rect 38 167 58 171
rect 65 167 77 171
rect 1 162 5 167
rect 20 162 24 167
rect 46 162 50 167
rect 84 162 88 171
rect -45 156 -30 162
rect -16 156 -9 162
rect -89 152 -85 156
rect -59 152 -55 156
rect 9 152 13 156
rect 28 152 32 156
rect 54 152 58 156
rect 73 152 77 156
rect -89 150 43 152
rect -89 146 -83 150
rect -79 146 -49 150
rect -45 146 15 150
rect 19 146 43 150
rect -89 144 43 146
rect 52 150 87 152
rect 52 146 60 150
rect 64 146 87 150
rect 52 144 87 146
rect -69 137 -15 141
rect -65 132 21 134
rect -65 128 -49 132
rect -45 128 14 132
rect 18 128 21 132
rect -65 126 21 128
rect 29 132 88 134
rect 29 128 61 132
rect 65 128 88 132
rect 29 126 88 128
rect -59 123 -55 126
rect -19 123 -15 126
rect 8 123 12 126
rect 28 123 32 126
rect 46 123 50 126
rect -45 115 -29 123
rect 54 123 58 126
rect 73 123 77 126
rect -29 112 -25 115
rect -9 112 -5 115
rect 19 112 23 115
rect 38 112 42 115
rect 65 112 69 115
rect 84 112 94 115
rect -29 108 12 112
rect 19 108 31 112
rect 38 108 58 112
rect 65 108 77 112
rect -9 103 -5 108
rect 19 103 23 108
rect 46 103 50 108
rect 84 103 88 112
rect -45 97 -29 103
rect -59 93 -55 97
rect 8 93 12 97
rect 28 93 32 97
rect 54 93 58 97
rect 73 93 77 97
rect -62 91 43 93
rect -62 87 -49 91
rect -45 87 13 91
rect 17 87 43 91
rect -62 85 43 87
rect 52 91 87 93
rect 52 87 59 91
rect 63 87 87 91
rect 52 85 87 87
rect -97 78 -5 82
rect -97 70 -92 74
rect -84 73 21 75
rect -84 69 -49 73
rect -45 69 15 73
rect 19 69 21 73
rect -84 67 21 69
rect 29 73 88 75
rect 29 69 61 73
rect 65 69 88 73
rect 29 67 88 69
rect -84 64 -80 67
rect -59 64 -55 67
rect -29 64 -25 67
rect 9 64 13 67
rect 28 64 32 67
rect 46 64 50 67
rect -45 56 -39 64
rect -25 56 -9 64
rect 54 64 58 67
rect 73 64 77 67
rect -68 51 -64 56
rect -39 53 -35 56
rect 1 53 5 56
rect 20 53 24 56
rect 38 53 42 56
rect 65 53 69 56
rect 84 53 94 56
rect -97 47 -83 51
rect -76 47 -64 51
rect -39 49 13 53
rect 20 49 31 53
rect 38 49 58 53
rect 65 49 77 53
rect -76 44 -72 47
rect 1 44 5 49
rect 20 44 24 49
rect 46 44 50 49
rect 84 44 88 53
rect -84 34 -80 38
rect -68 34 -64 38
rect -45 38 -39 44
rect -25 38 -9 44
rect -59 34 -55 38
rect 9 34 13 38
rect 28 34 32 38
rect 54 34 58 38
rect 73 34 77 38
rect -97 32 43 34
rect -97 28 -49 32
rect -45 28 15 32
rect 19 28 43 32
rect -97 26 43 28
rect 52 32 87 34
rect 52 28 60 32
rect 64 28 87 32
rect 52 26 87 28
rect -62 19 41 23
rect -97 13 21 15
rect -97 9 -49 13
rect -45 9 14 13
rect 18 9 21 13
rect -97 7 21 9
rect 29 13 88 15
rect 29 9 61 13
rect 65 9 88 13
rect 29 7 88 9
rect -83 4 -79 7
rect -59 4 -55 7
rect -29 4 -25 7
rect 8 4 12 7
rect 28 4 32 7
rect 46 4 50 7
rect -45 -4 -39 4
rect -25 -4 -19 4
rect 54 4 58 7
rect 73 4 77 7
rect -72 -7 -68 -4
rect -39 -7 -35 -4
rect -9 -7 -5 -4
rect 19 -7 23 -4
rect 38 -7 42 -4
rect 65 -7 69 -4
rect 84 -7 94 -4
rect -87 -11 -79 -7
rect -39 -11 12 -7
rect 19 -11 31 -7
rect 38 -11 58 -7
rect 65 -11 77 -7
rect -72 -16 -68 -12
rect -9 -16 -5 -11
rect 19 -16 23 -11
rect 46 -16 50 -11
rect 84 -16 88 -7
rect -45 -22 -39 -16
rect -25 -22 -19 -16
rect -83 -26 -79 -22
rect -59 -26 -55 -22
rect 8 -26 12 -22
rect 28 -26 32 -22
rect 54 -26 58 -22
rect 73 -26 77 -22
rect -97 -28 43 -26
rect -97 -32 -49 -28
rect -45 -32 13 -28
rect 17 -32 43 -28
rect -97 -34 43 -32
rect 52 -28 87 -26
rect 52 -32 59 -28
rect 63 -32 87 -28
rect 52 -34 87 -32
<< m2contact >>
rect 21 422 29 430
rect -74 403 -69 408
rect 65 399 70 404
rect 43 381 52 389
rect -74 373 -69 378
rect 21 363 29 371
rect 65 340 70 345
rect 43 322 52 330
rect 21 303 29 311
rect -74 284 -69 289
rect 65 280 70 285
rect 43 262 52 270
rect -74 254 -69 259
rect 21 244 29 252
rect 65 221 70 226
rect 43 203 52 211
rect 21 185 29 193
rect -74 166 -69 171
rect 65 162 70 167
rect 43 144 52 152
rect -74 136 -69 141
rect 21 126 29 134
rect 65 103 70 108
rect 43 85 52 93
rect 21 67 29 75
rect -64 47 -59 52
rect 65 44 70 49
rect 43 26 52 34
rect -67 18 -62 23
rect 21 7 29 15
rect -92 -11 -87 -6
rect -72 -12 -67 -7
rect 65 -16 70 -11
rect 43 -34 52 -26
<< metal2 >>
rect -74 378 -69 403
rect 21 371 29 422
rect 70 399 94 403
rect 21 311 29 363
rect -74 259 -69 284
rect 21 252 29 303
rect 21 193 29 244
rect -74 141 -69 166
rect 21 134 29 185
rect 21 75 29 126
rect -64 32 -59 47
rect -92 27 -59 32
rect -92 -6 -87 27
rect -67 -12 -62 18
rect 21 15 29 67
rect 43 330 52 381
rect 70 340 94 344
rect 43 270 52 322
rect 70 280 94 284
rect 43 211 52 262
rect 70 221 94 225
rect 43 152 52 203
rect 70 162 94 166
rect 43 93 52 144
rect 70 103 94 107
rect 43 34 52 85
rect 70 44 94 48
rect 43 -26 52 26
rect 70 -16 94 -12
<< labels >>
rlabel metal1 66 346 66 346 1 wl6
rlabel metal1 68 405 68 405 1 wl7
rlabel metal1 -96 406 -96 406 3 A
rlabel metal1 66 286 66 286 1 wl5
rlabel metal1 -96 287 -96 287 3 B
rlabel metal1 66 168 66 168 1 wl3
rlabel metal1 66 227 66 227 1 wl4
rlabel metal1 -96 169 -96 169 3 C
rlabel metal1 66 110 66 110 1 wl2
rlabel metal1 66 51 66 51 1 wl1
rlabel metal1 93 410 93 410 7 Nwl7
rlabel metal1 91 350 91 350 7 Nwl6
rlabel metal1 91 290 91 290 7 Nwl5
rlabel metal1 91 232 91 232 7 Nwl4
rlabel metal1 91 172 91 172 7 Nwl3
rlabel metal1 90 113 90 113 7 Nwl2
rlabel metal1 90 54 90 54 7 Nwl1
rlabel metal1 -58 11 -58 11 1 Vdd
rlabel metal1 -58 -30 -58 -30 1 Gnd
rlabel metal1 66 -9 66 -9 1 wl0
rlabel metal1 91 -5 91 -5 7 Nwl0
rlabel metal1 -94 72 -94 72 3 clear_r
rlabel metal1 -93 49 -93 49 3 calc_hist_r
<< end >>
