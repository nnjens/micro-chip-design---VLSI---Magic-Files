magic
tech scmos
timestamp 1480993349
<< polysilicon >>
rect 1184 469 1189 473
<< polycontact >>
rect 1189 468 1194 474
<< metal1 >>
rect 1709 1985 1865 1986
rect 243 1983 1865 1985
rect 243 1973 340 1983
rect 350 1974 1713 1983
rect 1722 1974 1865 1983
rect 350 1973 1865 1974
rect 368 1972 370 1973
rect 247 1669 378 1679
rect 391 1678 639 1679
rect 391 1669 992 1678
rect 14 1253 25 1260
rect 14 1226 19 1234
rect 22 1212 30 1218
rect 14 1106 19 1118
rect 361 1075 369 1092
rect 13 990 18 1002
rect 8 900 13 904
rect 21 877 22 881
rect 1174 481 1203 489
rect 1189 456 1194 468
rect 1194 435 1195 437
rect 791 419 795 429
rect 843 418 847 430
rect 895 418 899 430
rect 1188 429 1195 435
rect 926 419 934 423
rect 947 418 951 428
rect 999 418 1003 428
rect 1051 418 1055 428
rect 1103 418 1107 428
rect 1155 419 1159 429
rect 757 397 775 405
rect 935 398 1011 407
rect 1365 405 1370 409
rect 939 346 958 355
rect 968 346 993 355
rect 938 320 958 324
rect 1156 322 1173 326
rect 755 272 773 280
rect 924 278 1000 287
rect 937 219 958 228
rect 968 219 991 228
rect 1153 202 1170 206
rect 936 196 958 200
rect 934 169 1010 178
rect 752 154 770 162
rect 935 102 957 109
rect 967 102 969 109
rect 932 78 958 82
<< m2contact >>
rect 14 877 21 884
rect 1187 435 1194 444
rect 926 410 934 419
rect 958 346 968 355
rect 958 219 968 228
rect 957 102 967 111
<< metal2 >>
rect 8 932 16 933
rect 8 925 29 932
rect 22 884 29 925
rect 21 877 29 884
rect 1142 435 1187 443
rect 925 410 926 418
rect 934 410 968 418
rect 958 355 968 410
rect 958 228 968 346
rect 958 111 968 219
rect 967 103 968 111
<< m123contact >>
rect 340 1972 350 1983
rect 1713 1974 1722 1983
rect 378 1669 391 1679
rect 1712 1671 1721 1680
rect 369 1369 384 1377
rect 1708 1367 1722 1377
rect 13 1234 19 1241
rect 361 1092 369 1097
rect 1712 1069 1725 1078
rect 1368 457 1373 462
rect 764 370 770 377
rect 942 372 947 377
rect 981 373 986 378
rect 1160 374 1165 379
rect 764 247 769 253
rect 942 248 947 253
rect 981 253 986 258
rect 1160 254 1165 259
rect 764 129 769 135
rect 942 130 947 135
<< m234contact >>
rect 1 925 8 932
<< metal4 >>
rect 349 1972 350 1980
<< m345contact >>
rect 350 1972 359 1981
rect 1722 1974 1731 1983
rect 1712 1680 1721 1689
rect 367 1669 378 1679
rect 1708 1377 1722 1387
rect 369 1361 385 1369
rect 13 1227 19 1234
rect 369 1091 380 1097
rect 1709 1078 1721 1087
rect 158 768 167 775
rect 135 673 144 679
rect 13 604 25 616
rect 1368 462 1373 467
rect 942 377 947 382
rect 1160 379 1165 384
rect 758 370 764 377
rect 972 373 981 378
rect 1160 259 1165 264
rect 942 253 947 258
rect 972 253 981 258
rect 759 247 764 253
rect 136 206 147 220
rect 942 135 947 140
rect 759 129 764 135
<< metal5 >>
rect 349 1972 350 1980
rect 378 1669 383 1679
rect 370 1383 383 1669
rect 369 1377 383 1383
rect 369 1369 384 1377
rect 369 1321 383 1361
rect 15 1234 67 1236
rect 19 1227 67 1234
rect 15 1226 67 1227
rect 369 1097 384 1321
rect 380 1091 384 1097
rect 204 925 205 932
rect 167 768 169 775
rect 14 144 25 604
rect 135 258 144 673
rect 160 379 169 768
rect 194 688 205 925
rect 195 394 205 688
rect 369 664 384 1091
rect 942 382 952 620
rect 947 377 952 382
rect 942 258 952 377
rect 1160 384 1170 622
rect 1165 379 1170 384
rect 947 253 952 258
rect 1160 264 1170 379
rect 1165 259 1170 264
rect 942 140 952 253
rect 1160 251 1170 259
<< m456contact >>
rect 8 925 16 933
<< m6contact >>
rect 359 1972 370 1984
rect 1731 1974 1748 1983
rect 1696 1689 1721 1698
rect 356 1669 367 1679
rect 1696 1387 1722 1397
rect 194 925 204 933
rect 1696 1087 1721 1096
rect 369 618 410 664
rect 942 620 952 668
rect 1159 622 1170 677
rect 195 385 205 394
rect 160 370 169 379
rect 750 370 758 378
rect 973 378 981 386
rect 134 248 144 258
rect 1368 467 1376 475
rect 751 247 759 255
rect 972 258 980 266
rect 125 206 136 220
rect 14 132 25 144
rect 751 129 759 137
<< metal6 >>
rect 1705 1985 1722 1986
rect 358 1972 359 1980
rect 359 1687 370 1972
rect 1696 1983 1749 1985
rect 1696 1974 1731 1983
rect 1748 1974 1749 1983
rect 1696 1973 1749 1974
rect 1696 1698 1722 1973
rect 1721 1689 1722 1698
rect 356 1679 391 1687
rect 367 1669 391 1679
rect 1696 1397 1722 1689
rect 1696 1096 1722 1387
rect 1721 1087 1722 1096
rect 1696 1078 1722 1087
rect 1696 1069 1725 1078
rect 1696 1052 1722 1069
rect 16 925 194 933
rect 204 925 207 933
rect 369 664 942 665
rect 368 620 369 643
rect 410 620 942 664
rect 952 622 1159 665
rect 1696 665 1721 1052
rect 1170 622 1721 665
rect 952 620 1721 622
rect 410 619 1721 620
rect 410 618 1595 619
rect 1368 475 1377 618
rect 1695 516 1721 619
rect 1695 514 1720 516
rect 1376 467 1377 475
rect 405 395 986 396
rect 195 394 986 395
rect 205 386 986 394
rect 205 385 776 386
rect 160 379 759 380
rect 169 378 759 379
rect 169 370 750 378
rect 758 370 759 378
rect 108 266 980 274
rect 108 264 972 266
rect 108 220 123 264
rect 144 255 760 258
rect 144 248 751 255
rect 759 248 760 255
rect 108 206 125 220
rect 136 206 146 220
rect 108 205 146 206
rect 25 141 161 142
rect 25 137 759 141
rect 25 132 751 137
rect 14 131 751 132
use FF  FF_1
timestamp 1480480681
transform -1 0 909 0 -1 321
box -36 -84 140 28
use FF  FF_4
timestamp 1480480681
transform -1 0 1126 0 -1 323
box -36 -84 140 28
use FF  FF_0
timestamp 1480480681
transform -1 0 1334 0 -1 406
box -36 -84 140 28
use FF  FF_2
timestamp 1480480681
transform -1 0 908 0 -1 197
box -36 -84 140 28
use FF  FF_5
timestamp 1480480681
transform -1 0 1126 0 -1 203
box -36 -84 140 28
use FF  FF_3
timestamp 1480480681
transform -1 0 908 0 -1 79
box -36 -84 140 28
use d_m_mux_f  d_m_mux_f_0
timestamp 1480988083
transform 1 0 12 0 1 521
box -12 -521 2159 1532
<< labels >>
rlabel metal1 792 421 792 421 1 out_hist7
rlabel metal1 844 421 844 421 1 out_hist6
rlabel metal1 897 421 897 421 1 out_hist5
rlabel metal1 949 421 949 421 1 out_hist4
rlabel metal1 1002 421 1002 421 1 out_hist3
rlabel metal1 1053 421 1053 421 1 out_hist2
rlabel metal1 1105 421 1105 421 1 out_hist1
rlabel metal1 1156 421 1156 421 1 out_hist0
rlabel metal6 1715 540 1715 540 1 clk_top
rlabel metal1 956 322 956 322 1 input2
rlabel metal1 955 199 955 199 1 input1
rlabel metal1 952 80 952 80 1 input0
rlabel metal1 1172 324 1172 324 1 calc_hist
rlabel metal1 1166 204 1166 204 1 clear
rlabel polysilicon 1185 470 1185 470 1 out_valid
rlabel metal2 960 304 960 304 1 Gnd
rlabel metal1 765 276 765 276 1 Vdd
rlabel metal1 1367 407 1367 407 1 read_out
<< end >>
