magic
tech scmos
timestamp 1481052353
<< nwell >>
rect -50 -59 465 31
rect -50 -62 452 -59
<< pwell >>
rect 452 -62 465 -59
rect -50 -119 465 -62
<< ntransistor >>
rect -35 -78 -33 -73
rect -19 -103 -17 -68
rect -3 -103 -1 -68
rect 5 -103 7 -68
rect 13 -103 15 -68
rect 21 -103 23 -68
rect 29 -103 31 -68
rect 37 -103 39 -68
rect 45 -103 47 -68
rect 61 -103 63 -68
rect 69 -103 71 -68
rect 77 -103 79 -68
rect 85 -103 87 -68
rect 93 -103 95 -68
rect 101 -103 103 -68
rect 109 -103 111 -68
rect 117 -103 119 -68
rect 125 -103 127 -68
rect 133 -103 135 -68
rect 141 -103 143 -68
rect 149 -103 151 -68
rect 157 -103 159 -68
rect 165 -103 167 -68
rect 173 -103 175 -68
rect 181 -103 183 -68
rect 189 -103 191 -68
rect 197 -103 199 -68
rect 205 -103 207 -68
rect 213 -103 215 -68
rect 221 -103 223 -68
rect 229 -103 231 -68
rect 237 -103 239 -68
rect 245 -103 247 -68
rect 253 -103 255 -68
rect 261 -103 263 -68
rect 269 -103 271 -68
rect 277 -103 279 -68
rect 285 -103 287 -68
rect 293 -103 295 -68
rect 301 -103 303 -68
rect 309 -103 311 -68
rect 317 -103 319 -68
rect 325 -103 327 -68
rect 333 -103 335 -68
rect 341 -103 343 -68
rect 349 -103 351 -68
rect 357 -103 359 -68
rect 365 -103 367 -68
rect 373 -103 375 -68
rect 381 -103 383 -68
rect 389 -103 391 -68
rect 397 -103 399 -68
rect 405 -103 407 -68
rect 413 -103 415 -68
rect 421 -103 423 -68
rect 429 -103 431 -68
rect 437 -103 439 -68
rect 445 -103 447 -68
<< ptransistor >>
rect -35 -52 -33 -42
rect -19 -52 -17 18
rect -3 -52 -1 18
rect 5 -52 7 18
rect 13 -52 15 18
rect 21 -52 23 18
rect 29 -52 31 18
rect 37 -52 39 18
rect 45 -52 47 18
rect 61 -52 63 18
rect 69 -52 71 18
rect 77 -52 79 18
rect 85 -52 87 18
rect 93 -52 95 18
rect 101 -52 103 18
rect 109 -52 111 18
rect 117 -52 119 18
rect 125 -52 127 18
rect 133 -52 135 18
rect 141 -52 143 18
rect 149 -52 151 18
rect 157 -52 159 18
rect 165 -52 167 18
rect 173 -52 175 18
rect 181 -52 183 18
rect 189 -52 191 18
rect 197 -52 199 18
rect 205 -52 207 18
rect 213 -52 215 18
rect 221 -52 223 18
rect 229 -52 231 18
rect 237 -52 239 18
rect 245 -52 247 18
rect 253 -52 255 18
rect 261 -52 263 18
rect 269 -52 271 18
rect 277 -52 279 18
rect 285 -52 287 18
rect 293 -52 295 18
rect 301 -52 303 18
rect 309 -52 311 18
rect 317 -52 319 18
rect 325 -52 327 18
rect 333 -52 335 18
rect 341 -52 343 18
rect 349 -52 351 18
rect 357 -52 359 18
rect 365 -52 367 18
rect 373 -52 375 18
rect 381 -52 383 18
rect 389 -52 391 18
rect 397 -52 399 18
rect 405 -52 407 18
rect 413 -52 415 18
rect 421 -52 423 18
rect 429 -52 431 18
rect 437 -52 439 18
rect 445 -52 447 18
<< ndiffusion >>
rect -36 -78 -35 -73
rect -33 -78 -32 -73
rect -20 -103 -19 -68
rect -17 -103 -16 -68
rect -4 -103 -3 -68
rect -1 -103 5 -68
rect 7 -103 13 -68
rect 15 -103 21 -68
rect 23 -103 29 -68
rect 31 -103 37 -68
rect 39 -103 45 -68
rect 47 -103 48 -68
rect 60 -103 61 -68
rect 63 -103 69 -68
rect 71 -103 77 -68
rect 79 -103 85 -68
rect 87 -103 93 -68
rect 95 -103 101 -68
rect 103 -103 109 -68
rect 111 -103 117 -68
rect 119 -103 125 -68
rect 127 -103 133 -68
rect 135 -103 141 -68
rect 143 -103 149 -68
rect 151 -103 157 -68
rect 159 -103 165 -68
rect 167 -103 173 -68
rect 175 -103 181 -68
rect 183 -103 189 -68
rect 191 -103 197 -68
rect 199 -103 205 -68
rect 207 -103 213 -68
rect 215 -103 221 -68
rect 223 -103 229 -68
rect 231 -103 237 -68
rect 239 -103 245 -68
rect 247 -103 253 -68
rect 255 -103 261 -68
rect 263 -103 269 -68
rect 271 -103 277 -68
rect 279 -103 285 -68
rect 287 -103 293 -68
rect 295 -103 301 -68
rect 303 -103 309 -68
rect 311 -103 317 -68
rect 319 -103 325 -68
rect 327 -103 333 -68
rect 335 -103 341 -68
rect 343 -103 349 -68
rect 351 -103 357 -68
rect 359 -103 365 -68
rect 367 -103 373 -68
rect 375 -103 381 -68
rect 383 -103 389 -68
rect 391 -103 397 -68
rect 399 -103 405 -68
rect 407 -103 413 -68
rect 415 -103 421 -68
rect 423 -103 429 -68
rect 431 -103 437 -68
rect 439 -103 445 -68
rect 447 -103 448 -68
<< pdiffusion >>
rect -36 -52 -35 -42
rect -33 -52 -32 -42
rect -20 -52 -19 18
rect -17 -52 -16 18
rect -4 -52 -3 18
rect -1 -52 0 18
rect 4 -52 5 18
rect 7 -52 8 18
rect 12 -52 13 18
rect 15 -52 16 18
rect 20 -52 21 18
rect 23 -52 24 18
rect 28 -52 29 18
rect 31 -52 32 18
rect 36 -52 37 18
rect 39 -52 40 18
rect 44 -52 45 18
rect 47 -52 48 18
rect 60 -52 61 18
rect 63 -52 64 18
rect 68 -52 69 18
rect 71 -52 72 18
rect 76 -52 77 18
rect 79 -52 80 18
rect 84 -52 85 18
rect 87 -52 88 18
rect 92 -52 93 18
rect 95 -52 96 18
rect 100 -52 101 18
rect 103 -52 104 18
rect 108 -52 109 18
rect 111 -52 112 18
rect 116 -52 117 18
rect 119 -52 120 18
rect 124 -52 125 18
rect 127 -52 128 18
rect 132 -52 133 18
rect 135 -52 136 18
rect 140 -52 141 18
rect 143 -52 144 18
rect 148 -52 149 18
rect 151 -52 152 18
rect 156 -52 157 18
rect 159 -52 160 18
rect 164 -52 165 18
rect 167 -52 168 18
rect 172 -52 173 18
rect 175 -52 176 18
rect 180 -52 181 18
rect 183 -52 184 18
rect 188 -52 189 18
rect 191 -52 192 18
rect 196 -52 197 18
rect 199 -52 200 18
rect 204 -52 205 18
rect 207 -52 208 18
rect 212 -52 213 18
rect 215 -52 216 18
rect 220 -52 221 18
rect 223 -52 224 18
rect 228 -52 229 18
rect 231 -52 232 18
rect 236 -52 237 18
rect 239 -52 240 18
rect 244 -52 245 18
rect 247 -52 248 18
rect 252 -52 253 18
rect 255 -52 256 18
rect 260 -52 261 18
rect 263 -52 264 18
rect 268 -52 269 18
rect 271 -52 272 18
rect 276 -52 277 18
rect 279 -52 280 18
rect 284 -52 285 18
rect 287 -52 288 18
rect 292 -52 293 18
rect 295 -52 296 18
rect 300 -52 301 18
rect 303 -52 304 18
rect 308 -52 309 18
rect 311 -52 312 18
rect 316 -52 317 18
rect 319 -52 320 18
rect 324 -52 325 18
rect 327 -52 328 18
rect 332 -52 333 18
rect 335 -52 336 18
rect 340 -52 341 18
rect 343 -52 344 18
rect 348 -52 349 18
rect 351 -52 352 18
rect 356 -52 357 18
rect 359 -52 360 18
rect 364 -52 365 18
rect 367 -52 368 18
rect 372 -52 373 18
rect 375 -52 376 18
rect 380 -52 381 18
rect 383 -52 384 18
rect 388 -52 389 18
rect 391 -52 392 18
rect 396 -52 397 18
rect 399 -52 400 18
rect 404 -52 405 18
rect 407 -52 408 18
rect 412 -52 413 18
rect 415 -52 416 18
rect 420 -52 421 18
rect 423 -52 424 18
rect 428 -52 429 18
rect 431 -52 432 18
rect 436 -52 437 18
rect 439 -52 440 18
rect 444 -52 445 18
rect 447 -52 448 18
<< ndcontact >>
rect -40 -78 -36 -73
rect -32 -78 -28 -73
rect -24 -103 -20 -68
rect -16 -103 -12 -68
rect -8 -103 -4 -68
rect 48 -103 52 -68
rect 56 -103 60 -68
rect 448 -103 452 -68
<< pdcontact >>
rect -40 -52 -36 -42
rect -32 -52 -28 -42
rect -24 -52 -20 18
rect -16 -52 -12 18
rect -8 -52 -4 18
rect 0 -52 4 18
rect 8 -52 12 18
rect 16 -52 20 18
rect 24 -52 28 18
rect 32 -52 36 18
rect 40 -52 44 18
rect 48 -52 52 18
rect 56 -52 60 18
rect 64 -52 68 18
rect 72 -52 76 18
rect 80 -52 84 18
rect 88 -52 92 18
rect 96 -52 100 18
rect 104 -52 108 18
rect 112 -52 116 18
rect 120 -52 124 18
rect 128 -52 132 18
rect 136 -52 140 18
rect 144 -52 148 18
rect 152 -52 156 18
rect 160 -52 164 18
rect 168 -52 172 18
rect 176 -52 180 18
rect 184 -52 188 18
rect 192 -52 196 18
rect 200 -52 204 18
rect 208 -52 212 18
rect 216 -52 220 18
rect 224 -52 228 18
rect 232 -52 236 18
rect 240 -52 244 18
rect 248 -52 252 18
rect 256 -52 260 18
rect 264 -52 268 18
rect 272 -52 276 18
rect 280 -52 284 18
rect 288 -52 292 18
rect 296 -52 300 18
rect 304 -52 308 18
rect 312 -52 316 18
rect 320 -52 324 18
rect 328 -52 332 18
rect 336 -52 340 18
rect 344 -52 348 18
rect 352 -52 356 18
rect 360 -52 364 18
rect 368 -52 372 18
rect 376 -52 380 18
rect 384 -52 388 18
rect 392 -52 396 18
rect 400 -52 404 18
rect 408 -52 412 18
rect 416 -52 420 18
rect 424 -52 428 18
rect 432 -52 436 18
rect 440 -52 444 18
rect 448 -52 452 18
<< psubstratepcontact >>
rect -40 -115 452 -110
<< nsubstratencontact >>
rect -41 22 461 27
<< polysilicon >>
rect -19 18 -17 21
rect -3 18 -1 21
rect 5 18 7 21
rect 13 18 15 21
rect 21 18 23 21
rect 29 18 31 21
rect 37 18 39 21
rect 45 18 47 21
rect 61 18 63 21
rect 69 18 71 21
rect 77 18 79 21
rect 85 18 87 21
rect 93 18 95 21
rect 101 18 103 21
rect 109 18 111 21
rect 117 18 119 21
rect 125 18 127 21
rect 133 18 135 21
rect 141 18 143 21
rect 149 18 151 21
rect 157 18 159 21
rect 165 18 167 21
rect 173 18 175 21
rect 181 18 183 21
rect 189 18 191 21
rect 197 18 199 21
rect 205 18 207 21
rect 213 18 215 21
rect 221 18 223 21
rect 229 18 231 21
rect 237 18 239 21
rect 245 18 247 21
rect 253 18 255 21
rect 261 18 263 21
rect 269 18 271 21
rect 277 18 279 21
rect 285 18 287 21
rect 293 18 295 21
rect 301 18 303 21
rect 309 18 311 21
rect 317 18 319 21
rect 325 18 327 21
rect 333 18 335 21
rect 341 18 343 21
rect 349 18 351 21
rect 357 18 359 21
rect 365 18 367 21
rect 373 18 375 21
rect 381 18 383 21
rect 389 18 391 21
rect 397 18 399 21
rect 405 18 407 21
rect 413 18 415 21
rect 421 18 423 21
rect 429 18 431 21
rect 437 18 439 21
rect 445 18 447 21
rect -35 -42 -33 -39
rect -35 -73 -33 -52
rect -19 -68 -17 -52
rect -3 -56 -1 -52
rect 5 -56 7 -52
rect 13 -56 15 -52
rect 21 -56 23 -52
rect 29 -56 31 -52
rect 37 -56 39 -52
rect 45 -56 47 -52
rect -3 -63 47 -56
rect 61 -57 63 -52
rect 69 -57 71 -52
rect 77 -57 79 -52
rect 85 -57 87 -52
rect 93 -57 95 -52
rect 101 -57 103 -52
rect 109 -57 111 -52
rect 117 -57 119 -52
rect 125 -57 127 -52
rect 133 -57 135 -52
rect 141 -57 143 -52
rect 149 -57 151 -52
rect 157 -57 159 -52
rect 165 -57 167 -52
rect 173 -57 175 -52
rect 181 -57 183 -52
rect 189 -57 191 -52
rect 197 -57 199 -52
rect 205 -57 207 -52
rect 213 -57 215 -52
rect 221 -57 223 -52
rect 229 -57 231 -52
rect 237 -57 239 -52
rect 245 -57 247 -52
rect 253 -57 255 -52
rect 261 -57 263 -52
rect 269 -57 271 -52
rect 277 -57 279 -52
rect 285 -57 287 -52
rect 293 -57 295 -52
rect 301 -57 303 -52
rect 309 -57 311 -52
rect 317 -57 319 -52
rect 325 -57 327 -52
rect 333 -57 335 -52
rect 341 -57 343 -52
rect 349 -57 351 -52
rect 357 -57 359 -52
rect 365 -57 367 -52
rect 373 -57 375 -52
rect 381 -57 383 -52
rect 389 -57 391 -52
rect 397 -57 399 -52
rect 405 -57 407 -52
rect 413 -57 415 -52
rect 421 -57 423 -52
rect 429 -57 431 -52
rect 437 -57 439 -52
rect 445 -57 447 -52
rect -3 -68 -1 -63
rect 5 -68 7 -63
rect 13 -68 15 -63
rect 21 -68 23 -63
rect 29 -68 31 -63
rect 37 -68 39 -63
rect 45 -68 47 -63
rect 61 -64 447 -57
rect 61 -68 63 -64
rect 69 -68 71 -64
rect 77 -68 79 -64
rect 85 -68 87 -64
rect 93 -68 95 -64
rect 101 -68 103 -64
rect 109 -68 111 -64
rect 117 -68 119 -64
rect 125 -68 127 -64
rect 133 -68 135 -64
rect 141 -68 143 -64
rect 149 -68 151 -64
rect 157 -68 159 -64
rect 165 -68 167 -64
rect 173 -68 175 -64
rect 181 -68 183 -64
rect 189 -68 191 -64
rect 197 -68 199 -64
rect 205 -68 207 -64
rect 213 -68 215 -64
rect 221 -68 223 -64
rect 229 -68 231 -64
rect 237 -68 239 -64
rect 245 -68 247 -64
rect 253 -68 255 -64
rect 261 -68 263 -64
rect 269 -68 271 -64
rect 277 -68 279 -64
rect 285 -68 287 -64
rect 293 -68 295 -64
rect 301 -68 303 -64
rect 309 -68 311 -64
rect 317 -68 319 -64
rect 325 -68 327 -64
rect 333 -68 335 -64
rect 341 -68 343 -64
rect 349 -68 351 -64
rect 357 -68 359 -64
rect 365 -68 367 -64
rect 373 -68 375 -64
rect 381 -68 383 -64
rect 389 -68 391 -64
rect 397 -68 399 -64
rect 405 -68 407 -64
rect 413 -68 415 -64
rect 421 -68 423 -64
rect 429 -68 431 -64
rect 437 -68 439 -64
rect 445 -68 447 -64
rect -35 -81 -33 -78
rect -19 -106 -17 -103
rect -3 -106 -1 -103
rect 5 -106 7 -103
rect 13 -106 15 -103
rect 21 -106 23 -103
rect 29 -106 31 -103
rect 37 -106 39 -103
rect 45 -106 47 -103
rect 61 -106 63 -103
rect 69 -106 71 -103
rect 77 -106 79 -103
rect 85 -106 87 -103
rect 93 -106 95 -103
rect 101 -106 103 -103
rect 109 -106 111 -103
rect 117 -106 119 -103
rect 125 -106 127 -103
rect 133 -106 135 -103
rect 141 -106 143 -103
rect 149 -106 151 -103
rect 157 -106 159 -103
rect 165 -106 167 -103
rect 173 -106 175 -103
rect 181 -106 183 -103
rect 189 -106 191 -103
rect 197 -106 199 -103
rect 205 -106 207 -103
rect 213 -106 215 -103
rect 221 -106 223 -103
rect 229 -106 231 -103
rect 237 -106 239 -103
rect 245 -106 247 -103
rect 253 -106 255 -103
rect 261 -106 263 -103
rect 269 -106 271 -103
rect 277 -106 279 -103
rect 285 -106 287 -103
rect 293 -106 295 -103
rect 301 -106 303 -103
rect 309 -106 311 -103
rect 317 -106 319 -103
rect 325 -106 327 -103
rect 333 -106 335 -103
rect 341 -106 343 -103
rect 349 -106 351 -103
rect 357 -106 359 -103
rect 365 -106 367 -103
rect 373 -106 375 -103
rect 381 -106 383 -103
rect 389 -106 391 -103
rect 397 -106 399 -103
rect 405 -106 407 -103
rect 413 -106 415 -103
rect 421 -106 423 -103
rect 429 -106 431 -103
rect 437 -106 439 -103
rect 445 -106 447 -103
<< polycontact >>
rect -40 -63 -35 -58
rect -24 -62 -19 -57
rect -8 -62 -3 -57
rect 56 -62 61 -57
<< metal1 >>
rect -44 27 461 29
rect -44 22 -41 27
rect -44 21 461 22
rect -40 -42 -36 21
rect -24 18 -20 21
rect -8 18 -4 21
rect 8 18 12 21
rect 24 18 28 21
rect 40 18 44 21
rect 56 18 60 21
rect 72 18 76 21
rect 88 18 92 21
rect 104 18 108 21
rect 120 18 124 21
rect 136 18 140 21
rect 152 18 156 21
rect 168 18 172 21
rect 184 18 188 21
rect 200 18 204 21
rect 216 18 220 21
rect 232 18 236 21
rect 248 18 252 21
rect 264 18 268 21
rect 280 18 284 21
rect 296 18 300 21
rect 312 18 316 21
rect 328 18 332 21
rect 344 18 348 21
rect 360 18 364 21
rect 376 18 380 21
rect 392 18 396 21
rect 408 18 412 21
rect 424 18 428 21
rect 440 18 444 21
rect -32 -57 -28 -52
rect -16 -57 -12 -52
rect 0 -57 4 -52
rect 16 -57 20 -52
rect 32 -57 36 -52
rect 48 -57 52 -52
rect 64 -57 68 -52
rect 80 -57 84 -52
rect 96 -57 100 -52
rect 112 -57 116 -52
rect 128 -57 132 -52
rect 144 -57 148 -52
rect 160 -57 164 -52
rect 176 -57 180 -52
rect 192 -57 196 -52
rect 208 -57 212 -52
rect 224 -57 228 -52
rect 240 -57 244 -52
rect 256 -57 260 -52
rect 272 -57 276 -52
rect 288 -57 292 -52
rect 304 -57 308 -52
rect 320 -57 324 -52
rect 336 -57 340 -52
rect 352 -57 356 -52
rect 368 -57 372 -52
rect 384 -57 388 -52
rect 400 -57 404 -52
rect 416 -57 420 -52
rect 432 -57 436 -52
rect 448 -57 452 -52
rect -44 -63 -40 -58
rect -32 -62 -24 -57
rect -16 -62 -8 -57
rect 0 -62 56 -57
rect 64 -62 452 -57
rect -32 -73 -28 -62
rect -16 -68 -12 -62
rect 48 -68 52 -62
rect 448 -68 452 -62
rect -40 -109 -36 -78
rect -24 -109 -20 -103
rect -8 -109 -4 -103
rect 56 -109 60 -103
rect -50 -110 452 -109
rect -50 -115 -40 -110
rect -50 -117 452 -115
<< labels >>
rlabel metal1 450 -60 450 -60 1 out
rlabel metal1 -42 -61 -42 -61 1 in
rlabel nsubstratencontact -35 25 -35 25 1 Vdd
rlabel metal1 -44 -114 -44 -114 1 Gnd
<< end >>
