magic
tech scmos
timestamp 1480978990
<< nwell >>
rect 564 -323 569 -318
rect 640 -323 645 -318
rect 716 -325 721 -320
<< pwell >>
rect 810 -86 818 -79
rect 862 -86 870 -79
rect 914 -86 922 -79
rect 966 -86 974 -79
rect 1018 -86 1026 -79
rect 1070 -86 1078 -79
rect 1122 -86 1130 -79
rect 159 -381 164 -376
rect 235 -381 240 -376
rect 311 -381 316 -376
rect 387 -380 392 -375
rect 539 -380 544 -375
rect 615 -380 620 -375
<< polysilicon >>
rect 801 -52 1178 -48
rect 801 -56 804 -52
rect 853 -57 856 -52
rect 905 -57 908 -52
rect 957 -56 960 -52
rect 1009 -57 1012 -52
rect 1061 -56 1064 -52
rect 1114 -56 1117 -52
rect 1166 -54 1169 -52
<< metal1 >>
rect 229 1449 243 1459
rect 1110 1452 1123 1459
rect 236 1151 246 1157
rect 1110 1150 1122 1159
rect 246 847 261 856
rect 1108 849 1116 857
rect 4 731 16 739
rect 1 713 10 717
rect 10 690 15 698
rect 1 594 10 598
rect 238 548 258 554
rect 1109 550 1125 557
rect 1 476 9 480
rect -4 379 9 383
rect 3 356 14 360
rect 1087 155 1095 187
rect 1070 148 1095 155
rect 145 3 153 109
rect 763 27 774 28
rect 674 18 774 27
rect 762 -9 774 18
rect 142 -40 174 -36
rect 218 -40 251 -34
rect 295 -40 327 -34
rect 371 -40 403 -34
rect 446 -40 479 -35
rect 483 -37 487 -27
rect 559 -28 560 -25
rect 522 -40 555 -35
rect 559 -37 564 -28
rect 598 -39 631 -34
rect 675 -40 679 -35
rect 703 -37 707 -15
rect 728 -18 733 -10
rect 746 -16 774 -9
rect 862 16 893 26
rect 746 -18 773 -16
rect 862 -56 870 16
rect 986 -54 992 -7
rect 1038 -54 1043 -18
rect 1070 -60 1078 148
rect 1120 16 1161 26
rect 1121 -16 1130 16
rect 1211 -7 1220 27
rect 1163 -16 1221 -7
rect 1121 -22 1131 -16
rect 1091 -55 1095 -29
rect 1122 -56 1131 -22
rect 1142 -55 1147 -41
rect 1163 -64 1172 -16
rect 779 -102 783 -95
rect 831 -103 835 -96
rect 883 -103 887 -96
rect 935 -103 939 -96
rect 987 -103 991 -96
rect 1039 -103 1043 -96
rect 1091 -103 1095 -96
rect 1143 -102 1147 -95
rect 283 -350 286 -346
rect 142 -355 147 -352
rect 142 -359 173 -355
rect 142 -363 156 -359
rect 168 -360 173 -359
rect 168 -365 193 -360
rect 208 -364 212 -351
rect 218 -355 223 -350
rect 218 -359 248 -355
rect 218 -363 232 -359
rect 224 -364 232 -363
rect 243 -360 248 -359
rect 243 -364 269 -360
rect 283 -363 288 -350
rect 294 -355 299 -348
rect 294 -359 324 -355
rect 294 -363 309 -359
rect 320 -360 324 -359
rect 320 -364 345 -360
rect 357 -363 364 -349
rect 370 -354 375 -350
rect 370 -358 400 -354
rect 370 -362 384 -358
rect 395 -359 400 -358
rect 395 -363 421 -359
rect 435 -361 440 -349
rect 451 -353 476 -352
rect 446 -358 476 -353
rect 446 -360 460 -358
rect 452 -362 460 -360
rect 471 -363 497 -358
rect 508 -362 516 -345
rect 585 -346 589 -345
rect 522 -352 527 -349
rect 522 -358 551 -352
rect 522 -362 536 -358
rect 547 -363 573 -358
rect 584 -361 592 -346
rect 598 -352 603 -345
rect 662 -347 668 -346
rect 598 -358 628 -352
rect 598 -362 612 -358
rect 623 -363 649 -358
rect 660 -362 668 -347
rect 674 -352 679 -348
rect 674 -358 705 -352
rect 674 -362 689 -358
rect 403 -364 418 -363
rect 700 -364 726 -358
rect 737 -363 744 -345
<< m2contact >>
rect 179 -37 184 -29
rect 255 -39 260 -32
rect 933 -55 940 -49
rect 758 -86 766 -79
rect 810 -86 818 -79
rect 862 -86 870 -79
rect 914 -86 922 -79
rect 966 -86 974 -79
rect 1018 -86 1026 -79
rect 1070 -86 1078 -79
rect 1122 -86 1130 -79
rect 741 -98 747 -91
rect 799 -98 807 -91
rect 851 -98 859 -91
rect 903 -98 911 -91
rect 955 -98 963 -91
rect 1007 -98 1015 -91
rect 1059 -98 1067 -91
rect 1111 -98 1119 -91
rect 1163 -98 1171 -91
rect 184 -324 189 -319
rect 260 -326 265 -321
rect 336 -323 341 -318
rect 412 -325 417 -320
rect 488 -326 493 -321
rect 564 -323 569 -318
rect 640 -323 645 -318
rect 716 -325 721 -320
<< metal2 >>
rect 404 21 621 27
rect 126 -11 131 18
rect 255 12 392 18
rect 399 12 400 18
rect 126 -16 178 -11
rect 179 -29 183 -18
rect 255 -32 259 12
rect 404 8 410 21
rect 616 18 621 21
rect 331 3 410 8
rect 432 10 611 17
rect 616 14 664 18
rect 933 12 938 24
rect 933 10 940 12
rect 179 -44 183 -37
rect 255 -44 259 -39
rect 331 -43 336 3
rect 432 -1 438 10
rect 607 4 940 10
rect 407 -7 438 -1
rect 407 -47 412 -7
rect 674 -32 737 -27
rect 732 -39 737 -32
rect 933 -49 940 4
rect 766 -86 810 -79
rect 818 -86 862 -79
rect 870 -86 914 -79
rect 922 -86 966 -79
rect 974 -86 1018 -79
rect 1026 -86 1070 -79
rect 1078 -86 1122 -79
rect 747 -98 799 -91
rect 807 -98 851 -91
rect 859 -98 903 -91
rect 911 -98 955 -91
rect 963 -98 1007 -91
rect 1015 -98 1059 -91
rect 1067 -98 1111 -91
rect 1119 -92 1125 -91
rect 1119 -98 1163 -92
rect 565 -318 569 -313
rect 189 -324 190 -322
rect 185 -360 190 -324
rect 341 -323 342 -319
rect 261 -360 265 -326
rect 177 -365 190 -360
rect 253 -364 265 -360
rect 337 -361 342 -323
rect 417 -325 418 -321
rect 413 -359 418 -325
rect 493 -326 494 -322
rect 489 -359 494 -326
rect 565 -359 569 -323
rect 329 -365 344 -361
rect 405 -364 420 -359
rect 481 -363 494 -359
rect 557 -364 569 -359
rect 641 -360 645 -323
rect 633 -364 645 -360
rect 717 -361 721 -325
rect 709 -365 721 -361
rect 348 -435 353 -428
<< m3contact >>
rect 288 1451 295 1461
rect 388 1450 398 1460
rect 491 1451 501 1461
rect 594 1451 604 1461
rect 698 1451 708 1461
rect 800 1451 810 1461
rect 902 1452 913 1462
rect 1006 1452 1016 1462
rect 1201 10 1208 18
rect 1468 8 1476 18
rect 1739 7 1747 17
rect 2008 11 2015 18
rect 196 -438 201 -433
rect 272 -441 278 -432
rect 348 -446 354 -435
rect 424 -440 429 -429
rect 499 -440 506 -432
rect 576 -438 581 -429
rect 652 -442 657 -428
rect 729 -440 735 -430
<< m123contact >>
rect -12 378 -4 383
rect 483 -27 488 -22
rect 560 -28 565 -23
rect 635 -36 641 -31
rect 711 -48 716 -43
rect 984 -7 993 0
rect 1035 -18 1045 -11
rect 1089 -29 1098 -22
rect 1140 -41 1150 -34
rect 778 -56 784 -51
rect 830 -56 836 -51
rect 883 -56 889 -51
rect 159 -381 164 -376
rect 235 -381 240 -376
rect 311 -381 316 -376
rect 387 -380 392 -375
rect 463 -380 468 -375
rect 539 -380 544 -375
rect 615 -380 620 -375
rect 692 -380 697 -375
<< metal3 >>
rect -12 77 -4 378
rect -12 71 78 77
rect 71 16 78 71
rect 71 7 135 16
rect 2008 18 2015 21
rect 23 -514 31 -25
rect 35 -503 43 -25
rect 48 -491 56 -23
rect 60 -480 68 -22
rect 72 -467 80 -24
rect 84 -455 92 -23
rect 97 -444 105 -21
rect 110 -433 118 -19
rect 124 -375 135 7
rect 1202 1 1208 10
rect 1068 0 1208 1
rect 483 -7 984 0
rect 993 -7 1208 0
rect 1740 17 1746 18
rect 483 -22 488 -7
rect 1468 -11 1476 8
rect 559 -18 1035 -11
rect 1045 -18 1476 -11
rect 559 -23 565 -18
rect 1740 -22 1746 7
rect 559 -26 560 -23
rect 635 -29 1089 -22
rect 1098 -29 1746 -22
rect 635 -31 641 -29
rect 2008 -34 2015 11
rect 748 -41 1140 -34
rect 1150 -41 2015 -34
rect 748 -43 755 -41
rect 716 -47 755 -43
rect 716 -48 748 -47
rect 124 -376 387 -375
rect 124 -381 159 -376
rect 164 -381 235 -376
rect 240 -381 311 -376
rect 316 -380 387 -376
rect 392 -380 463 -375
rect 468 -380 539 -375
rect 544 -380 615 -375
rect 620 -380 692 -375
rect 316 -381 550 -380
rect 652 -428 657 -426
rect 576 -429 581 -428
rect 110 -438 196 -433
rect 110 -440 201 -438
rect 272 -444 277 -441
rect 97 -451 277 -444
rect 348 -455 353 -446
rect 84 -462 353 -455
rect 286 -463 353 -462
rect 424 -466 429 -440
rect 371 -467 429 -466
rect 72 -475 429 -467
rect 499 -432 506 -429
rect 72 -476 80 -475
rect 499 -480 506 -440
rect 60 -487 506 -480
rect 576 -491 581 -438
rect 48 -498 581 -491
rect 652 -503 657 -442
rect 35 -510 657 -503
rect 727 -440 729 -431
rect 727 -514 734 -440
rect 23 -521 734 -514
<< m234contact >>
rect 392 12 399 18
rect 664 14 670 20
rect 178 -18 185 -11
<< m4contact >>
rect 1006 1462 1016 1472
rect 281 1450 288 1460
rect 378 1450 388 1460
rect 481 1451 491 1461
rect 584 1451 594 1461
rect 688 1451 698 1461
rect 790 1451 800 1461
rect 893 1451 902 1461
rect 23 -25 31 -17
rect 35 -25 43 -17
rect 48 -23 56 -15
rect 60 -22 68 -14
rect 72 -24 80 -16
rect 84 -23 92 -15
rect 97 -21 105 -13
rect 110 -19 118 -11
rect 778 -51 784 -46
rect 830 -51 836 -46
rect 883 -51 889 -46
<< metal4 >>
rect 126 1531 263 1532
rect 124 1526 1017 1531
rect 124 1518 132 1526
rect 261 1525 1017 1526
rect 125 1449 131 1518
rect 138 1516 903 1520
rect 137 1514 903 1516
rect 125 1424 132 1449
rect 126 892 132 1424
rect 22 883 132 892
rect 22 798 31 883
rect 126 882 132 883
rect 137 878 143 1514
rect 36 875 143 878
rect 23 -17 31 798
rect 35 869 143 875
rect 148 1504 803 1510
rect 35 798 44 869
rect 49 864 126 865
rect 148 864 154 1504
rect 49 856 154 864
rect 49 834 56 856
rect 137 855 154 856
rect 158 1499 687 1500
rect 158 1494 700 1499
rect 158 850 164 1494
rect 170 1489 595 1490
rect 35 -17 43 798
rect 48 -15 56 834
rect 60 841 164 850
rect 60 -14 68 841
rect 158 840 164 841
rect 169 1484 595 1489
rect 169 836 175 1484
rect 72 827 175 836
rect 179 1474 491 1480
rect 72 -16 80 827
rect 179 823 185 1474
rect 84 822 166 823
rect 176 822 185 823
rect 84 814 185 822
rect 189 1464 389 1470
rect 84 -15 92 814
rect 189 808 195 1464
rect 378 1460 389 1464
rect 200 1451 281 1460
rect 200 1449 209 1451
rect 288 1451 296 1460
rect 388 1450 389 1460
rect 480 1461 491 1474
rect 480 1458 481 1461
rect 583 1461 594 1484
rect 583 1458 584 1461
rect 688 1461 699 1494
rect 789 1462 802 1504
rect 790 1461 801 1462
rect 800 1456 801 1461
rect 893 1461 902 1514
rect 1006 1472 1016 1525
rect 199 1398 209 1449
rect 199 1394 210 1398
rect 200 1196 210 1394
rect 97 799 195 808
rect 199 1191 210 1196
rect 97 -13 105 799
rect 199 794 209 1191
rect 110 785 209 794
rect 111 410 119 785
rect 110 404 119 410
rect 110 -11 118 404
rect 853 20 859 21
rect 670 14 860 20
rect 392 3 399 12
rect 392 -3 837 3
rect 778 -11 784 -10
rect 185 -17 786 -11
rect 778 -46 784 -17
rect 831 -46 836 -3
rect 853 -41 859 14
rect 853 -46 889 -41
rect 853 -47 883 -46
rect 778 -55 784 -51
rect 831 -54 836 -51
rect 883 -54 887 -51
use d_m_mux  d_m_mux_0
timestamp 1480978990
transform 1 0 36 0 1 259
box -36 -259 2123 1201
use fadder8  fadder8_0
timestamp 1480976721
transform 0 1 724 -1 0 -8
box -14 -584 349 27
use AND  AND_0
timestamp 1480867771
transform 0 1 789 -1 0 -68
box -15 -31 33 19
use AND  AND_1
timestamp 1480867771
transform 0 1 841 -1 0 -68
box -15 -31 33 19
use AND  AND_2
timestamp 1480867771
transform 0 1 893 -1 0 -68
box -15 -31 33 19
use AND  AND_3
timestamp 1480867771
transform 0 1 945 -1 0 -68
box -15 -31 33 19
use AND  AND_4
timestamp 1480867771
transform 0 1 997 -1 0 -68
box -15 -31 33 19
use AND  AND_5
timestamp 1480867771
transform 0 1 1049 -1 0 -68
box -15 -31 33 19
use AND  AND_6
timestamp 1480867771
transform 0 1 1101 -1 0 -68
box -15 -31 33 19
use AND  AND_7
timestamp 1480867771
transform 0 1 1153 -1 0 -68
box -15 -31 33 19
use mux21  mux21_0
timestamp 1480737015
transform 0 1 165 -1 0 -403
box -41 -18 31 47
use mux21  mux21_1
timestamp 1480737015
transform 0 1 241 -1 0 -403
box -41 -18 31 47
use mux21  mux21_2
timestamp 1480737015
transform 0 1 317 -1 0 -403
box -41 -18 31 47
use mux21  mux21_3
timestamp 1480737015
transform 0 1 393 -1 0 -402
box -41 -18 31 47
use mux21  mux21_4
timestamp 1480737015
transform 0 1 469 -1 0 -402
box -41 -18 31 47
use mux21  mux21_5
timestamp 1480737015
transform 0 1 545 -1 0 -402
box -41 -18 31 47
use mux21  mux21_6
timestamp 1480737015
transform 0 1 621 -1 0 -402
box -41 -18 31 47
use mux21  mux21_7
timestamp 1480737015
transform 0 1 698 -1 0 -402
box -41 -18 31 47
<< labels >>
rlabel metal3 -9 375 -9 375 3 clear_r
rlabel metal1 6 357 6 358 1 calc_hist_r
rlabel metal1 4 478 4 478 1 input0_r
rlabel metal1 2 596 2 596 1 input1_r
rlabel metal1 2 715 2 715 1 input2_r
rlabel metal1 11 735 11 736 1 Vdd
rlabel metal1 12 694 12 694 1 Gnd
rlabel polysilicon 1176 -51 1176 -51 1 read_out_r
rlabel metal1 781 -100 781 -100 1 out_hist7
rlabel metal1 833 -101 833 -101 1 out_hist6
rlabel metal1 885 -101 885 -101 1 out_hist5
rlabel metal1 937 -100 937 -100 1 out_hist4
rlabel metal1 989 -100 989 -100 1 out_hist3
rlabel metal1 1041 -100 1041 -100 1 out_hist2
rlabel metal1 1093 -100 1093 -100 1 out_hist1
rlabel metal1 1145 -100 1145 -100 1 out_hist0
rlabel metal1 239 1153 239 1153 1 clk1
rlabel metal1 234 1450 234 1450 1 clk0
rlabel metal1 253 851 253 851 1 clk2
rlabel metal1 240 549 240 549 1 clk3
rlabel metal1 1114 1456 1114 1456 1 clk4
rlabel metal1 1114 1157 1114 1157 1 clk5
rlabel metal1 1112 856 1112 856 1 clk6
rlabel metal1 1112 555 1112 555 1 clk7
<< end >>
