magic
tech scmos
timestamp 1480562330
<< nwell >>
rect -56 -501 -24 -451
rect 25 -501 79 -451
rect 128 -501 182 -451
rect 231 -501 285 -451
rect 334 -501 388 -451
rect 437 -501 491 -451
rect 540 -501 594 -451
rect 643 -501 697 -451
rect 665 -506 697 -501
rect 746 -506 777 -451
<< pwell >>
rect -24 -501 25 -451
rect 79 -501 128 -451
rect 182 -501 231 -451
rect 285 -501 334 -451
rect 388 -501 437 -451
rect 491 -501 540 -451
rect 594 -501 643 -451
rect 697 -506 746 -451
<< ntransistor >>
rect -11 -486 -7 -484
rect 9 -486 13 -484
rect 92 -486 96 -484
rect 112 -486 116 -484
rect 195 -486 199 -484
rect 215 -486 219 -484
rect 298 -486 302 -484
rect 318 -486 322 -484
rect 401 -486 405 -484
rect 421 -486 425 -484
rect 504 -486 508 -484
rect 524 -486 528 -484
rect 607 -486 611 -484
rect 627 -486 631 -484
rect 710 -486 714 -484
rect 730 -486 734 -484
<< ptransistor >>
rect -43 -486 -37 -484
rect 36 -486 42 -484
rect 60 -486 66 -484
rect 139 -486 145 -484
rect 163 -486 169 -484
rect 242 -486 248 -484
rect 266 -486 272 -484
rect 345 -486 351 -484
rect 369 -486 375 -484
rect 448 -486 454 -484
rect 472 -486 478 -484
rect 551 -486 557 -484
rect 575 -486 581 -484
rect 654 -486 660 -484
rect 678 -486 684 -484
rect 757 -486 763 -484
<< ndiffusion >>
rect -11 -484 -7 -483
rect 9 -484 13 -483
rect -11 -487 -7 -486
rect 9 -487 13 -486
rect 92 -484 96 -483
rect 112 -484 116 -483
rect 92 -487 96 -486
rect 112 -487 116 -486
rect 195 -484 199 -483
rect 215 -484 219 -483
rect 195 -487 199 -486
rect 215 -487 219 -486
rect 298 -484 302 -483
rect 318 -484 322 -483
rect 298 -487 302 -486
rect 318 -487 322 -486
rect 401 -484 405 -483
rect 421 -484 425 -483
rect 401 -487 405 -486
rect 421 -487 425 -486
rect 504 -484 508 -483
rect 524 -484 528 -483
rect 504 -487 508 -486
rect 524 -487 528 -486
rect 607 -484 611 -483
rect 627 -484 631 -483
rect 607 -487 611 -486
rect 627 -487 631 -486
rect 710 -484 714 -483
rect 730 -484 734 -483
rect 710 -487 714 -486
rect 730 -487 734 -486
<< pdiffusion >>
rect -43 -484 -37 -483
rect -43 -487 -37 -486
rect 36 -484 42 -483
rect 60 -484 66 -483
rect 36 -487 42 -486
rect 60 -487 66 -486
rect 139 -484 145 -483
rect 163 -484 169 -483
rect 139 -487 145 -486
rect 163 -487 169 -486
rect 242 -484 248 -483
rect 266 -484 272 -483
rect 242 -487 248 -486
rect 266 -487 272 -486
rect 345 -484 351 -483
rect 369 -484 375 -483
rect 345 -487 351 -486
rect 369 -487 375 -486
rect 448 -484 454 -483
rect 472 -484 478 -483
rect 448 -487 454 -486
rect 472 -487 478 -486
rect 551 -484 557 -483
rect 575 -484 581 -483
rect 551 -487 557 -486
rect 575 -487 581 -486
rect 654 -484 660 -483
rect 678 -484 684 -483
rect 654 -487 660 -486
rect 678 -487 684 -486
rect 757 -484 763 -483
rect 757 -487 763 -486
<< polysilicon >>
rect -46 -486 -43 -484
rect -37 -486 -34 -484
rect -14 -486 -11 -484
rect -7 -486 -4 -484
rect 6 -486 9 -484
rect 13 -486 16 -484
rect 33 -486 36 -484
rect 42 -486 45 -484
rect 57 -486 60 -484
rect 66 -486 69 -484
rect 89 -486 92 -484
rect 96 -486 99 -484
rect 109 -486 112 -484
rect 116 -486 119 -484
rect 136 -486 139 -484
rect 145 -486 148 -484
rect 160 -486 163 -484
rect 169 -486 172 -484
rect 192 -486 195 -484
rect 199 -486 202 -484
rect 212 -486 215 -484
rect 219 -486 222 -484
rect 239 -486 242 -484
rect 248 -486 251 -484
rect 263 -486 266 -484
rect 272 -486 275 -484
rect 295 -486 298 -484
rect 302 -486 305 -484
rect 315 -486 318 -484
rect 322 -486 325 -484
rect 342 -486 345 -484
rect 351 -486 354 -484
rect 366 -486 369 -484
rect 375 -486 378 -484
rect 398 -486 401 -484
rect 405 -486 408 -484
rect 418 -486 421 -484
rect 425 -486 428 -484
rect 445 -486 448 -484
rect 454 -486 457 -484
rect 469 -486 472 -484
rect 478 -486 481 -484
rect 501 -486 504 -484
rect 508 -486 511 -484
rect 521 -486 524 -484
rect 528 -486 531 -484
rect 548 -486 551 -484
rect 557 -486 560 -484
rect 572 -486 575 -484
rect 581 -486 584 -484
rect 604 -486 607 -484
rect 611 -486 614 -484
rect 624 -486 627 -484
rect 631 -486 634 -484
rect 651 -486 654 -484
rect 660 -486 663 -484
rect 675 -486 678 -484
rect 684 -486 687 -484
rect 707 -486 710 -484
rect 714 -486 717 -484
rect 727 -486 730 -484
rect 734 -486 737 -484
rect 754 -486 757 -484
rect 763 -486 766 -484
<< polycontact >>
rect -34 -487 -30 -483
rect -18 -487 -14 -483
rect 16 -487 20 -483
rect 29 -487 33 -483
rect 69 -487 73 -483
rect 85 -487 89 -483
rect 119 -487 123 -483
rect 132 -487 136 -483
rect 172 -487 176 -483
rect 188 -487 192 -483
rect 222 -487 226 -483
rect 235 -487 239 -483
rect 275 -487 279 -483
rect 291 -487 295 -483
rect 325 -487 329 -483
rect 338 -487 342 -483
rect 378 -487 382 -483
rect 394 -487 398 -483
rect 428 -487 432 -483
rect 441 -487 445 -483
rect 481 -487 485 -483
rect 497 -487 501 -483
rect 531 -487 535 -483
rect 544 -487 548 -483
rect 584 -487 588 -483
rect 600 -487 604 -483
rect 634 -487 638 -483
rect 647 -487 651 -483
rect 687 -487 691 -483
rect 703 -487 707 -483
rect 737 -487 741 -483
rect 750 -487 754 -483
<< metal1 >>
rect -25 -448 700 -441
rect -55 -503 -47 -457
rect -34 -483 -30 -465
rect -25 -470 -21 -448
rect -27 -476 -21 -470
rect -27 -502 -23 -476
rect -18 -483 -14 -474
rect -3 -501 5 -457
rect 16 -483 20 -460
rect 29 -483 33 -469
rect 47 -501 55 -457
rect 69 -483 73 -465
rect 78 -468 82 -448
rect 76 -473 82 -468
rect 76 -501 80 -473
rect 85 -483 89 -474
rect 100 -501 108 -457
rect 119 -483 123 -460
rect 132 -483 136 -469
rect 150 -501 158 -457
rect 172 -483 176 -465
rect 181 -468 185 -448
rect 179 -475 185 -468
rect 179 -501 183 -475
rect 188 -483 192 -474
rect 203 -501 211 -457
rect 222 -483 226 -460
rect 235 -483 239 -469
rect 253 -501 261 -457
rect 275 -483 279 -465
rect 284 -469 288 -448
rect 282 -474 288 -469
rect 282 -501 286 -474
rect 291 -483 295 -474
rect 306 -501 314 -457
rect 325 -483 329 -460
rect 338 -483 342 -469
rect 356 -501 364 -457
rect 378 -483 382 -465
rect 387 -468 391 -448
rect 385 -474 391 -468
rect 385 -501 389 -474
rect 394 -483 398 -474
rect 409 -501 417 -457
rect 428 -483 432 -460
rect 441 -483 445 -469
rect 459 -501 467 -457
rect 481 -483 485 -465
rect 490 -470 494 -448
rect 488 -474 494 -470
rect 488 -502 492 -474
rect 497 -483 501 -474
rect 512 -501 520 -457
rect 531 -483 535 -460
rect 544 -483 548 -469
rect 562 -501 570 -457
rect 584 -483 588 -465
rect 593 -469 597 -448
rect 591 -477 597 -469
rect 591 -501 595 -477
rect 600 -483 604 -474
rect 615 -501 623 -457
rect 634 -483 638 -460
rect 647 -483 651 -469
rect -55 -506 -48 -503
rect 665 -506 673 -454
rect 687 -483 691 -465
rect 696 -469 700 -448
rect 694 -474 700 -469
rect 694 -501 698 -474
rect 703 -483 707 -474
rect 718 -506 726 -457
rect 737 -483 741 -460
rect 750 -483 754 -463
rect 768 -503 776 -454
rect 24 -720 28 -716
rect 127 -720 131 -717
rect 230 -720 234 -716
rect 333 -720 337 -716
rect 436 -720 440 -716
rect 539 -720 543 -716
rect 642 -720 646 -716
rect 745 -720 749 -716
<< m2contact >>
rect 24 -501 29 -496
rect 127 -501 132 -496
rect 230 -501 235 -496
rect 333 -501 338 -496
rect 436 -501 441 -496
rect 539 -501 544 -496
rect 642 -501 647 -496
rect 745 -501 750 -496
rect -3 -685 5 -677
rect 100 -685 108 -677
rect 203 -685 211 -677
rect 306 -685 314 -677
rect 409 -685 417 -677
rect 512 -685 520 -677
rect 615 -685 623 -677
rect 718 -685 726 -677
<< pdm12contact >>
rect -43 -483 -37 -478
rect -43 -492 -37 -487
rect 36 -483 42 -478
rect 36 -492 42 -487
rect 60 -483 66 -478
rect 60 -492 66 -487
rect 139 -483 145 -478
rect 139 -492 145 -487
rect 163 -483 169 -478
rect 163 -492 169 -487
rect 242 -483 248 -478
rect 242 -492 248 -487
rect 266 -483 272 -478
rect 266 -492 272 -487
rect 345 -483 351 -478
rect 345 -492 351 -487
rect 369 -483 375 -478
rect 369 -492 375 -487
rect 448 -483 454 -478
rect 448 -492 454 -487
rect 472 -483 478 -478
rect 472 -492 478 -487
rect 551 -483 557 -478
rect 551 -492 557 -487
rect 575 -483 581 -478
rect 575 -492 581 -487
rect 654 -483 660 -478
rect 654 -492 660 -487
rect 678 -483 684 -478
rect 678 -492 684 -487
rect 757 -483 763 -478
rect 757 -492 763 -487
<< ndm12contact >>
rect -11 -483 -6 -478
rect -11 -492 -6 -487
rect 8 -483 13 -478
rect 8 -492 13 -487
rect 92 -483 97 -478
rect 92 -492 97 -487
rect 111 -483 116 -478
rect 111 -492 116 -487
rect 195 -483 200 -478
rect 195 -492 200 -487
rect 214 -483 219 -478
rect 214 -492 219 -487
rect 298 -483 303 -478
rect 298 -492 303 -487
rect 317 -483 322 -478
rect 317 -492 322 -487
rect 401 -483 406 -478
rect 401 -492 406 -487
rect 420 -483 425 -478
rect 420 -492 425 -487
rect 504 -483 509 -478
rect 504 -492 509 -487
rect 523 -483 528 -478
rect 523 -492 528 -487
rect 607 -483 612 -478
rect 607 -492 612 -487
rect 626 -483 631 -478
rect 626 -492 631 -487
rect 710 -483 715 -478
rect 710 -492 715 -487
rect 729 -483 734 -478
rect 729 -492 734 -487
<< metal2 >>
rect 23 -478 27 -464
rect 126 -478 130 -464
rect 229 -478 233 -464
rect 332 -478 336 -464
rect 435 -478 439 -464
rect 538 -478 542 -464
rect 641 -478 645 -464
rect 744 -478 748 -464
rect -37 -482 -27 -478
rect -22 -482 -11 -478
rect 13 -482 36 -478
rect 66 -482 76 -478
rect 81 -482 92 -478
rect 116 -482 139 -478
rect 169 -482 179 -478
rect 184 -482 195 -478
rect 219 -482 242 -478
rect 272 -482 282 -478
rect 287 -482 298 -478
rect 322 -482 345 -478
rect 375 -482 385 -478
rect 390 -482 401 -478
rect 425 -482 448 -478
rect 478 -482 488 -478
rect 493 -482 504 -478
rect 528 -482 551 -478
rect 581 -482 591 -478
rect 596 -482 607 -478
rect 631 -482 654 -478
rect 684 -482 694 -478
rect 699 -482 710 -478
rect 734 -482 757 -478
rect -37 -492 -11 -488
rect 13 -492 36 -488
rect 66 -492 92 -488
rect 116 -492 139 -488
rect 169 -492 195 -488
rect 219 -492 242 -488
rect 272 -492 298 -488
rect 322 -492 345 -488
rect 375 -492 401 -488
rect 425 -492 448 -488
rect 478 -492 504 -488
rect 528 -492 551 -488
rect 581 -492 607 -488
rect 631 -492 654 -488
rect 684 -492 710 -488
rect 734 -492 757 -488
rect -18 -496 -13 -492
rect 24 -496 29 -492
rect -18 -501 24 -496
rect 85 -496 90 -492
rect 127 -496 132 -492
rect 85 -501 127 -496
rect 188 -496 193 -492
rect 230 -496 235 -492
rect 188 -501 230 -496
rect 291 -496 296 -492
rect 333 -496 338 -492
rect 291 -501 333 -496
rect 394 -496 399 -492
rect 436 -496 441 -492
rect 394 -501 436 -496
rect 497 -496 502 -492
rect 539 -496 544 -492
rect 497 -501 539 -496
rect 600 -496 605 -492
rect 642 -496 647 -492
rect 600 -501 642 -496
rect 703 -496 708 -492
rect 745 -496 750 -492
rect 703 -501 745 -496
rect 5 -685 100 -677
rect 108 -685 203 -677
rect 211 -685 306 -677
rect 314 -685 409 -677
rect 417 -685 512 -677
rect 520 -685 615 -677
rect 623 -685 718 -677
<< m3contact >>
rect -27 -483 -22 -478
rect 76 -483 81 -478
rect 179 -483 184 -478
rect 282 -483 287 -478
rect 385 -483 390 -478
rect 488 -483 493 -478
rect 591 -483 596 -478
rect 694 -483 699 -478
<< m123contact >>
rect -34 -465 -29 -460
rect 11 -465 16 -460
rect -18 -474 -13 -469
rect 69 -465 74 -460
rect 114 -465 119 -460
rect 33 -474 38 -469
rect 85 -474 90 -469
rect 172 -465 177 -460
rect 217 -465 222 -460
rect 136 -474 141 -469
rect 188 -474 193 -469
rect 275 -465 280 -460
rect 320 -465 325 -460
rect 239 -474 244 -469
rect 291 -474 296 -469
rect 378 -465 383 -460
rect 423 -465 428 -460
rect 342 -474 347 -469
rect 394 -474 399 -469
rect 481 -465 486 -460
rect 526 -465 531 -460
rect 445 -474 450 -469
rect 497 -474 502 -469
rect 584 -465 589 -460
rect 629 -465 634 -460
rect 548 -474 553 -469
rect 600 -474 605 -469
rect 687 -465 692 -460
rect 732 -465 737 -460
rect 651 -474 656 -469
rect 703 -474 708 -469
rect 754 -474 759 -469
rect 23 -716 28 -711
rect 126 -716 131 -711
rect 229 -716 234 -711
rect 332 -716 337 -711
rect 435 -716 440 -711
rect 538 -716 543 -711
rect 641 -716 646 -711
rect 744 -716 749 -711
<< metal3 >>
rect -29 -465 11 -460
rect 16 -465 69 -460
rect 74 -465 114 -460
rect 119 -465 172 -460
rect 177 -465 217 -460
rect 222 -465 275 -460
rect 280 -465 320 -460
rect 325 -465 378 -460
rect 383 -465 423 -460
rect 428 -465 481 -460
rect 486 -465 526 -460
rect 531 -465 584 -460
rect 589 -465 629 -460
rect 634 -465 687 -460
rect 692 -465 732 -460
rect -13 -474 33 -469
rect 38 -474 85 -469
rect 90 -474 136 -469
rect 141 -474 188 -469
rect 193 -474 239 -469
rect 244 -474 291 -469
rect 296 -474 342 -469
rect 347 -474 394 -469
rect 399 -474 445 -469
rect 450 -474 497 -469
rect 502 -474 548 -469
rect 553 -474 600 -469
rect 605 -474 651 -469
rect 656 -474 703 -469
rect 708 -474 754 -469
rect -27 -711 -23 -483
rect 76 -711 80 -483
rect 179 -711 183 -483
rect 282 -711 286 -483
rect 385 -711 389 -483
rect 488 -711 492 -483
rect 591 -711 595 -483
rect 694 -711 698 -483
rect -27 -716 23 -711
rect 76 -716 126 -711
rect 179 -716 229 -711
rect 282 -716 332 -711
rect 385 -716 435 -711
rect 488 -716 538 -711
rect 591 -716 641 -711
rect 694 -716 744 -711
use buffer2  buffer2_6
timestamp 1480552228
transform 0 1 -56 -1 0 -497
box 0 0 224 112
use buffer2  buffer2_5
timestamp 1480552228
transform 0 1 47 -1 0 -497
box 0 0 224 112
use buffer2  buffer2_4
timestamp 1480552228
transform 0 1 150 -1 0 -497
box 0 0 224 112
use buffer2  buffer2_3
timestamp 1480552228
transform 0 1 253 -1 0 -497
box 0 0 224 112
use buffer2  buffer2_2
timestamp 1480552228
transform 0 1 356 -1 0 -497
box 0 0 224 112
use buffer2  buffer2_1
timestamp 1480552228
transform 0 1 459 -1 0 -497
box 0 0 224 112
use buffer2  buffer2_0
timestamp 1480552228
transform 0 1 562 -1 0 -497
box 0 0 224 112
use buffer  buffer_0
timestamp 1480483750
transform 0 1 665 -1 0 -497
box 0 0 224 112
<< labels >>
rlabel metal1 644 -718 644 -718 1 q1
rlabel metal1 541 -718 541 -718 1 q2
rlabel metal1 438 -718 438 -718 1 q3
rlabel metal1 335 -719 335 -719 1 q4
rlabel metal1 232 -717 232 -717 1 q5
rlabel metal1 129 -719 129 -719 1 q6
rlabel metal1 26 -719 26 -719 1 q7
rlabel metal1 747 -719 747 -719 1 q0
rlabel metal1 772 -462 772 -462 7 Vdd
rlabel metal1 752 -465 752 -465 3 Nen
rlabel metal1 739 -461 739 -461 3 en
rlabel metal2 746 -465 746 -465 3 new0
rlabel metal2 643 -467 643 -467 3 new1
rlabel metal2 540 -467 540 -467 3 new2
rlabel metal2 436 -466 436 -466 3 new3
rlabel metal2 334 -467 334 -467 3 new4
rlabel metal2 231 -467 231 -467 3 new5
rlabel metal2 128 -467 128 -467 3 new6
rlabel metal2 25 -467 25 -467 3 new7
rlabel metal1 723 -467 723 -467 3 Gnd
rlabel metal1 697 -443 697 -443 5 clk
<< end >>
