magic
tech scmos
timestamp 1480820178
<< nwell >>
rect 216 29 222 31
<< metal1 >>
rect 259 1177 267 1185
rect 1139 1179 1147 1186
rect 321 902 325 905
rect 1295 902 1299 906
rect 1398 902 1402 906
rect 1501 903 1505 907
rect 1604 903 1608 907
rect 1707 903 1711 907
rect 1810 903 1814 908
rect 1913 903 1917 908
rect 424 899 428 901
rect 527 897 531 900
rect 630 898 634 901
rect 733 898 737 901
rect 836 899 840 902
rect 939 899 943 902
rect 1042 899 1046 901
rect 1192 898 1196 901
rect 265 878 271 884
rect 1138 878 1146 885
rect 321 601 325 606
rect 424 601 428 606
rect 527 599 531 604
rect 630 598 634 603
rect 733 598 737 605
rect 836 597 840 604
rect 939 597 943 604
rect 1042 597 1046 604
rect 1192 596 1196 603
rect 1295 597 1299 604
rect 1398 597 1402 604
rect 1501 601 1505 608
rect 1604 600 1608 607
rect 1707 600 1711 604
rect 1810 602 1814 607
rect 1913 601 1917 606
rect 267 576 274 582
rect 1138 576 1148 583
rect 39 458 43 466
rect 215 458 243 466
rect 213 444 222 448
rect 30 440 33 444
rect 201 440 209 444
rect 212 443 222 444
rect 212 440 216 443
rect 39 417 43 425
rect 214 417 224 425
rect 215 399 243 407
rect 213 385 222 389
rect 202 381 209 385
rect 212 384 222 385
rect 212 381 216 384
rect 216 339 244 347
rect 30 321 33 325
rect 201 321 209 325
rect 212 324 222 329
rect 212 321 216 324
rect 321 297 325 303
rect 424 298 428 304
rect 527 299 531 305
rect 630 299 634 305
rect 733 298 737 305
rect 836 296 840 303
rect 939 295 943 302
rect 1042 296 1046 303
rect 1192 296 1196 304
rect 1295 295 1299 303
rect 1398 295 1402 303
rect 1501 295 1505 303
rect 1604 296 1608 305
rect 1707 299 1711 308
rect 1810 299 1814 308
rect 1913 300 1917 309
rect 215 280 243 288
rect 265 275 272 281
rect 1139 276 1150 283
rect 213 266 222 270
rect 200 262 209 266
rect 212 265 222 266
rect 212 262 216 265
rect 214 221 242 229
rect 213 207 222 211
rect 30 203 33 207
rect 202 203 209 207
rect 212 206 222 207
rect 212 203 216 206
rect 214 169 242 170
rect 214 162 244 169
rect 213 148 222 153
rect 201 144 209 148
rect 212 144 216 148
rect 31 106 34 110
rect 213 103 244 111
rect 213 88 222 93
rect 31 83 34 87
rect 214 43 245 51
rect 216 29 222 34
rect 211 2 234 10
rect 224 -1 234 2
rect 293 -1 301 4
rect 320 -1 324 4
rect 224 -10 301 -1
rect 423 -2 427 3
rect 526 -2 530 3
rect 629 -1 633 4
rect 732 -2 736 2
rect 835 -1 839 3
rect 938 -1 942 3
rect 1041 -2 1045 2
rect 1191 1 1195 6
rect 1294 1 1298 6
rect 1397 0 1401 5
rect 1500 1 1504 6
rect 1603 0 1607 6
rect 1706 0 1710 6
rect 1809 1 1813 7
rect 1912 1 1916 7
<< m2contact >>
rect 294 461 302 468
rect 224 417 232 425
<< metal2 >>
rect 320 1184 324 1187
rect 423 1182 427 1187
rect 526 1184 530 1187
rect 629 1184 633 1187
rect 732 1184 736 1187
rect 835 1184 839 1187
rect 938 1184 942 1187
rect 1041 1184 1045 1187
rect 234 462 294 468
rect 234 425 242 462
rect 262 461 294 462
rect 232 417 242 425
<< m3contact >>
rect 222 434 227 439
rect 222 375 227 380
rect 222 315 227 320
rect 222 256 227 261
rect 222 197 227 202
rect 222 138 227 143
rect 222 79 227 84
rect 222 20 227 25
<< m123contact >>
rect 222 443 227 448
rect 222 384 227 389
rect 222 324 227 329
rect 222 265 227 270
rect 222 206 227 211
rect 222 148 227 153
rect 222 88 227 93
rect 222 29 227 34
<< metal3 >>
rect 1117 259 1131 264
<< m4contact >>
rect 246 1161 251 1166
rect 1184 1162 1190 1167
rect 255 1152 260 1157
rect 1174 1153 1180 1158
rect 278 860 283 865
rect 1164 861 1170 866
rect 273 851 278 856
rect 1144 852 1150 857
rect 283 558 288 563
rect 1143 559 1149 564
rect 294 549 299 554
rect 1132 550 1138 555
rect 227 443 232 448
rect 227 434 232 439
rect 227 384 232 389
rect 227 375 232 380
rect 227 324 232 329
rect 227 315 232 320
rect 227 265 232 270
rect 227 256 232 261
rect 284 258 289 263
rect 1111 259 1117 265
rect 249 249 255 254
rect 1122 249 1128 255
rect 227 206 232 211
rect 227 197 232 202
rect 227 148 232 153
rect 227 138 232 143
rect 227 88 232 93
rect 227 79 232 84
rect 227 29 232 34
rect 227 20 232 25
<< metal4 >>
rect 246 508 251 1161
rect 163 503 251 508
rect 163 25 168 503
rect 255 499 260 1152
rect 172 494 260 499
rect 264 860 278 865
rect 172 34 177 494
rect 264 490 269 860
rect 181 485 269 490
rect 1150 852 1159 857
rect 181 84 186 485
rect 273 481 278 851
rect 190 476 278 481
rect 190 93 195 476
rect 283 472 288 558
rect 200 467 288 472
rect 200 143 205 467
rect 294 463 299 549
rect 209 458 299 463
rect 209 153 214 458
rect 232 443 1128 448
rect 232 434 1117 439
rect 232 384 1102 389
rect 232 375 1092 380
rect 232 324 1082 329
rect 232 315 1072 320
rect 227 277 1061 283
rect 227 270 232 277
rect 236 267 1051 273
rect 236 261 241 267
rect 232 256 241 261
rect 249 211 255 249
rect 232 206 255 211
rect 284 202 289 258
rect 232 197 289 202
rect 1045 197 1051 267
rect 1055 207 1061 277
rect 1066 217 1072 315
rect 1076 227 1082 324
rect 1086 236 1092 375
rect 1096 245 1102 384
rect 1111 265 1117 434
rect 1122 255 1128 443
rect 1132 245 1138 550
rect 1096 240 1138 245
rect 1143 236 1149 559
rect 1086 231 1149 236
rect 1153 227 1159 852
rect 1076 221 1159 227
rect 1164 217 1170 861
rect 1066 211 1170 217
rect 1174 207 1180 1153
rect 1055 201 1180 207
rect 1184 197 1190 1162
rect 1045 191 1190 197
rect 209 148 227 153
rect 200 138 227 143
rect 190 88 227 93
rect 181 79 227 84
rect 172 29 227 34
rect 163 20 227 25
use decoder  decoder_0
timestamp 1480810385
transform 1 0 128 0 1 36
box -98 -35 94 431
use memory  memory_0
timestamp 1480631328
transform 1 0 241 0 1 905
box -9 -907 1704 282
<< labels >>
rlabel metal1 31 442 31 442 3 input2_r
rlabel metal1 31 323 31 323 3 input1_r
rlabel metal1 30 203 33 207 3 input0_r
rlabel metal1 32 108 32 108 3 clear_r
rlabel metal1 32 85 32 85 3 calc_hist_r
rlabel metal2 322 1186 322 1186 5 new7
rlabel metal2 424 1186 424 1186 5 new6
rlabel metal2 527 1186 527 1186 5 new5
rlabel metal2 630 1186 630 1186 5 new4
rlabel metal2 733 1186 733 1186 5 new3
rlabel metal2 836 1186 836 1186 5 new2
rlabel metal2 939 1186 939 1186 5 new1
rlabel metal2 1043 1186 1043 1186 5 new0
rlabel metal1 323 904 323 904 1 Q0_7
rlabel metal1 426 900 426 900 1 Q0_6
rlabel metal1 529 899 529 899 1 Q0_5
rlabel metal1 632 899 632 899 1 Q0_4
rlabel metal1 735 900 735 900 1 Q0_3
rlabel metal1 838 900 838 900 1 Q0_2
rlabel metal1 941 900 941 900 1 Q0_1
rlabel metal1 1044 900 1044 900 1 Q0_0
rlabel metal1 1194 900 1194 900 1 Q4_7
rlabel metal1 1297 905 1297 905 1 Q4_6
rlabel metal1 1400 904 1400 904 1 Q4_5
rlabel metal1 1503 905 1503 905 1 Q4_4
rlabel metal1 1606 905 1606 905 1 Q4_3
rlabel metal1 1709 905 1709 905 1 Q4_2
rlabel metal1 1812 905 1812 905 1 Q4_1
rlabel metal1 1915 905 1915 905 1 Q4_0
rlabel metal1 322 603 322 603 1 Q1_7
rlabel metal1 426 603 426 603 1 Q1_6
rlabel metal1 529 602 529 602 1 Q1_5
rlabel metal1 632 599 632 599 1 Q1_4
rlabel metal1 735 599 735 599 1 Q1_3
rlabel metal1 838 597 838 599 1 Q1_2
rlabel metal1 941 598 941 598 1 Q1_1
rlabel metal1 1044 598 1044 598 1 Q1_0
rlabel metal1 1194 598 1194 598 1 Q5_7
rlabel metal1 1297 599 1297 599 1 Q5_6
rlabel metal1 1399 599 1399 599 1 Q5_5
rlabel metal1 1503 602 1503 602 1 Q5_4
rlabel metal1 1605 603 1605 603 1 Q5_3
rlabel metal1 1709 602 1709 602 1 Q5_2
rlabel metal1 1812 604 1812 604 1 Q5_1
rlabel metal1 1915 604 1915 604 1 Q5_0
rlabel metal1 323 302 323 302 1 Q2_7
rlabel metal1 426 301 426 301 1 Q2_6
rlabel metal1 529 302 529 302 1 Q2_5
rlabel metal1 632 302 632 302 1 Q2_4
rlabel metal1 735 301 735 301 1 Q2_3
rlabel metal1 838 297 838 297 1 Q2_2
rlabel metal1 941 297 941 297 1 Q2_1
rlabel metal1 1044 297 1044 297 1 Q2_0
rlabel metal1 1194 297 1194 298 1 Q6_7
rlabel metal1 1297 296 1297 297 1 Q6_6
rlabel metal1 1400 296 1400 297 1 Q6_5
rlabel metal1 1503 296 1503 297 1 Q6_4
rlabel metal1 1606 297 1606 297 1 Q6_3
rlabel metal1 1709 301 1709 301 1 Q6_2
rlabel metal1 1813 301 1813 301 1 Q6_1
rlabel metal1 1915 302 1915 302 1 Q6_0
rlabel metal1 322 1 322 1 1 Q3_7
rlabel metal1 426 0 426 0 1 Q3_6
rlabel metal1 528 0 528 0 1 Q3_5
rlabel metal1 1193 2 1193 2 1 Q7_7
rlabel metal1 1296 2 1296 2 1 Q7_6
rlabel metal1 1399 1 1399 1 1 Q7_5
rlabel metal1 1502 2 1502 2 1 Q7_4
rlabel metal1 1605 2 1605 2 1 Q7_3
rlabel metal1 1707 2 1707 2 1 Q7_2
rlabel metal1 1914 2 1914 2 1 Q7_0
rlabel metal1 631 1 631 1 1 Q3_4
rlabel metal1 735 0 735 0 1 Q3_3
rlabel metal1 837 1 837 1 1 Q3_2
rlabel metal1 939 1 939 1 1 Q3_1
rlabel metal1 1043 -1 1043 -1 1 Q3_0
rlabel metal1 263 1181 263 1181 1 clk0
rlabel metal1 267 881 267 881 1 clk1
rlabel metal1 270 579 270 579 1 clk2
rlabel metal1 267 276 267 276 1 clk3
rlabel metal1 1141 282 1141 282 1 clk7
rlabel metal1 1141 582 1141 582 1 clk6
rlabel metal1 1140 884 1140 884 1 clk5
rlabel metal1 1141 1183 1141 1183 5 clk4
rlabel metal1 1811 2 1811 2 1 Q7_1
rlabel metal1 41 462 41 462 1 Vdd
rlabel metal1 40 421 40 421 1 Gnd
<< end >>
