magic
tech scmos
timestamp 1481054774
<< nwell >>
rect -1006 2433 -972 2472
rect -759 2433 -725 2472
rect -1006 2432 -977 2433
rect -759 2431 -728 2433
rect -1834 1898 -1799 1904
rect -1834 1870 -1793 1898
rect -1834 1732 -1799 1739
rect -1836 1731 -1799 1732
rect -1836 1705 -1795 1731
rect -1835 945 -1800 953
rect -1835 919 -1795 945
rect 1028 596 1069 622
rect 1034 589 1069 596
rect -2322 327 -2321 333
rect 191 -241 217 -236
rect 184 -276 217 -241
<< pwell >>
rect -1035 2433 -1006 2472
rect -788 2433 -759 2472
rect -1027 2432 -1006 2433
rect -780 2432 -759 2433
rect -1834 1849 -1793 1870
rect -1834 1841 -1799 1849
rect -1835 1684 -1795 1705
rect -1835 1676 -1799 1684
rect -1835 898 -1795 919
rect -1835 890 -1800 898
rect 1034 648 1069 651
rect 1028 622 1069 648
rect -2322 383 -2321 390
rect -1237 182 -1229 199
rect 217 -241 238 -236
rect 217 -276 246 -241
<< ntransistor >>
rect -1017 2459 -1012 2461
rect -770 2459 -765 2461
rect -1017 2443 -1012 2445
rect -770 2443 -765 2445
rect -1823 1859 -1821 1864
rect -1807 1859 -1805 1864
rect -1824 1694 -1822 1699
rect -1808 1694 -1806 1699
rect -1824 908 -1822 913
rect -1808 908 -1806 913
rect 1040 628 1042 633
rect 1056 628 1058 633
rect 223 -249 228 -247
rect 223 -265 228 -263
<< ptransistor >>
rect -1000 2459 -990 2461
rect -753 2459 -743 2461
rect -1000 2443 -990 2445
rect -753 2443 -743 2445
rect -1823 1876 -1821 1886
rect -1807 1876 -1805 1886
rect -1824 1711 -1822 1721
rect -1808 1711 -1806 1721
rect -1824 925 -1822 935
rect -1808 925 -1806 935
rect 1040 606 1042 616
rect 1056 606 1058 616
rect 201 -249 211 -247
rect 201 -265 211 -263
<< ndiffusion >>
rect -1017 2461 -1012 2462
rect -770 2461 -765 2462
rect -1017 2458 -1012 2459
rect -770 2458 -765 2459
rect -1017 2445 -1012 2446
rect -770 2445 -765 2446
rect -1017 2442 -1012 2443
rect -770 2442 -765 2443
rect -1824 1859 -1823 1864
rect -1821 1859 -1820 1864
rect -1808 1859 -1807 1864
rect -1805 1859 -1804 1864
rect -1825 1694 -1824 1699
rect -1822 1694 -1821 1699
rect -1809 1694 -1808 1699
rect -1806 1694 -1805 1699
rect -1825 908 -1824 913
rect -1822 908 -1821 913
rect -1809 908 -1808 913
rect -1806 908 -1805 913
rect 1039 628 1040 633
rect 1042 628 1043 633
rect 1055 628 1056 633
rect 1058 628 1059 633
rect 223 -247 228 -246
rect 223 -250 228 -249
rect 223 -263 228 -262
rect 223 -266 228 -265
<< pdiffusion >>
rect -1000 2461 -990 2462
rect -753 2461 -743 2462
rect -1000 2458 -990 2459
rect -753 2458 -743 2459
rect -1000 2445 -990 2446
rect -753 2445 -743 2446
rect -1000 2442 -990 2443
rect -753 2442 -743 2443
rect -1824 1876 -1823 1886
rect -1821 1876 -1820 1886
rect -1808 1876 -1807 1886
rect -1805 1876 -1804 1886
rect -1825 1711 -1824 1721
rect -1822 1711 -1821 1721
rect -1809 1711 -1808 1721
rect -1806 1711 -1805 1721
rect -1825 925 -1824 935
rect -1822 925 -1821 935
rect -1809 925 -1808 935
rect -1806 925 -1805 935
rect 1039 606 1040 616
rect 1042 606 1043 616
rect 1055 606 1056 616
rect 1058 606 1059 616
rect 201 -247 211 -246
rect 201 -250 211 -249
rect 201 -263 211 -262
rect 201 -266 211 -265
<< ndcontact >>
rect -1017 2462 -1012 2466
rect -770 2462 -765 2466
rect -1017 2454 -1012 2458
rect -770 2454 -765 2458
rect -1017 2446 -1012 2450
rect -770 2446 -765 2450
rect -1017 2438 -1012 2442
rect -770 2438 -765 2442
rect -1828 1859 -1824 1864
rect -1820 1859 -1816 1864
rect -1812 1859 -1808 1864
rect -1804 1859 -1800 1864
rect -1829 1694 -1825 1699
rect -1821 1694 -1817 1699
rect -1813 1694 -1809 1699
rect -1805 1694 -1801 1699
rect -1829 908 -1825 913
rect -1821 908 -1817 913
rect -1813 908 -1809 913
rect -1805 908 -1801 913
rect 1035 628 1039 633
rect 1043 628 1047 633
rect 1051 628 1055 633
rect 1059 628 1063 633
rect 223 -246 228 -242
rect 223 -254 228 -250
rect 223 -262 228 -258
rect 223 -270 228 -266
<< pdcontact >>
rect -1000 2462 -990 2466
rect -753 2462 -743 2466
rect -1000 2454 -990 2458
rect -753 2454 -743 2458
rect -1000 2446 -990 2450
rect -753 2446 -743 2450
rect -1000 2438 -990 2442
rect -753 2438 -743 2442
rect -1828 1876 -1824 1886
rect -1820 1876 -1816 1886
rect -1812 1876 -1808 1886
rect -1804 1876 -1800 1886
rect -1829 1711 -1825 1721
rect -1821 1711 -1817 1721
rect -1813 1711 -1809 1721
rect -1805 1711 -1801 1721
rect -1829 925 -1825 935
rect -1821 925 -1817 935
rect -1813 925 -1809 935
rect -1805 925 -1801 935
rect 1035 606 1039 616
rect 1043 606 1047 616
rect 1051 606 1055 616
rect 1059 606 1063 616
rect 201 -246 211 -242
rect 201 -254 211 -250
rect 201 -262 211 -258
rect 201 -270 211 -266
<< psubstratepcontact >>
rect 265 219 269 556
<< nsubstratencontact >>
rect 218 212 223 550
<< polysilicon >>
rect -1020 2459 -1017 2461
rect -1012 2459 -1000 2461
rect -990 2459 -987 2461
rect -773 2459 -770 2461
rect -765 2459 -753 2461
rect -743 2459 -740 2461
rect -1024 2443 -1017 2445
rect -1012 2443 -1000 2445
rect -990 2443 -983 2445
rect -777 2443 -770 2445
rect -765 2443 -753 2445
rect -743 2443 -736 2445
rect -1823 1886 -1821 1889
rect -1807 1886 -1805 1893
rect -1823 1864 -1821 1876
rect -1807 1864 -1805 1876
rect -1823 1856 -1821 1859
rect -1807 1852 -1805 1859
rect -1824 1721 -1822 1724
rect -1808 1721 -1806 1728
rect -1824 1699 -1822 1711
rect -1808 1699 -1806 1711
rect -1824 1691 -1822 1694
rect -1808 1687 -1806 1694
rect -1824 935 -1822 938
rect -1808 935 -1806 942
rect -1824 913 -1822 925
rect -1808 913 -1806 925
rect -1824 905 -1822 908
rect -1808 901 -1806 908
rect 1040 633 1042 640
rect 1056 633 1058 636
rect 1040 616 1042 628
rect 1056 616 1058 628
rect 1040 599 1042 606
rect 1056 603 1058 606
rect 194 -249 201 -247
rect 211 -249 223 -247
rect 228 -249 235 -247
rect 198 -265 201 -263
rect 211 -265 223 -263
rect 228 -265 231 -263
<< polycontact >>
rect -1009 2461 -1003 2466
rect -762 2461 -756 2466
rect -1008 2445 -1004 2449
rect -761 2445 -757 2449
rect -1828 1867 -1823 1873
rect -1811 1868 -1807 1872
rect -1829 1702 -1824 1708
rect -1812 1703 -1808 1707
rect -1829 916 -1824 922
rect -1812 917 -1808 921
rect 1042 620 1046 624
rect 1058 619 1063 625
rect 215 -253 219 -249
rect 214 -270 220 -265
<< metal1 >>
rect -1496 3041 -1442 3046
rect -1506 3019 -1442 3041
rect -1497 3014 -1442 3019
rect -1506 2982 -1442 3014
rect -1281 3041 -1227 3046
rect -1291 3019 -1227 3041
rect -1282 3014 -1227 3019
rect -1291 2982 -1227 3014
rect -1498 2962 -1450 2966
rect -1283 2962 -1235 2966
rect -1476 2960 -1463 2962
rect -1261 2960 -1245 2962
rect -1474 2959 -1463 2960
rect -1260 2959 -1245 2960
rect -1471 2946 -1463 2959
rect -1254 2945 -1245 2959
rect -1028 2567 -974 2572
rect -1038 2545 -974 2567
rect -1029 2540 -974 2545
rect -1038 2509 -974 2540
rect -781 2567 -727 2572
rect -791 2545 -727 2567
rect -782 2540 -727 2545
rect -791 2509 -727 2540
rect -563 2569 -509 2574
rect -573 2547 -509 2569
rect -564 2542 -509 2547
rect -573 2510 -509 2542
rect -289 2570 -235 2575
rect -299 2548 -235 2570
rect -290 2543 -235 2548
rect -299 2511 -235 2543
rect -1034 2485 -978 2491
rect -787 2485 -731 2491
rect -1030 2479 -982 2485
rect -783 2479 -735 2485
rect -1026 2475 -986 2479
rect -779 2475 -739 2479
rect -1020 2472 -992 2475
rect -773 2472 -745 2475
rect -1035 2466 -1027 2472
rect -1009 2466 -1003 2472
rect -980 2466 -972 2472
rect -1035 2462 -1017 2466
rect -1468 2449 -1463 2455
rect -1416 2442 -1408 2456
rect -1252 2445 -1244 2455
rect -1035 2450 -1027 2462
rect -990 2462 -972 2466
rect -1012 2454 -1000 2458
rect -1035 2446 -1017 2450
rect -1008 2449 -1004 2454
rect -980 2450 -972 2462
rect -1035 2437 -1027 2446
rect -990 2446 -972 2450
rect -1012 2439 -1000 2442
rect -1012 2438 -1008 2439
rect -1003 2438 -1000 2439
rect -980 2437 -972 2446
rect -788 2466 -780 2472
rect -762 2466 -756 2472
rect -733 2466 -725 2472
rect -788 2462 -770 2466
rect -788 2450 -780 2462
rect -743 2462 -725 2466
rect -765 2454 -753 2458
rect -788 2446 -770 2450
rect -761 2449 -757 2454
rect -733 2450 -725 2462
rect -788 2437 -780 2446
rect -743 2446 -725 2450
rect -765 2438 -753 2442
rect -1035 2426 -1027 2430
rect -733 2437 -725 2446
rect -788 2426 -780 2430
rect -1751 2379 -1527 2409
rect -1497 2379 -1301 2409
rect -1271 2379 -1061 2409
rect -1031 2379 -982 2409
rect -970 2379 -849 2409
rect -818 2379 -735 2409
rect -723 2379 -581 2409
rect -551 2379 -341 2409
rect -311 2379 321 2409
rect 351 2379 699 2409
rect 729 2379 939 2409
rect 969 2379 1009 2409
rect -2405 2052 -2341 2106
rect -2400 2051 -2341 2052
rect -2400 2042 -2378 2051
rect -2373 2042 -2341 2051
rect -2325 2089 -2323 2098
rect -2325 2081 -2305 2089
rect -2325 2050 -2323 2081
rect -1781 2015 -1751 2379
rect -1781 1906 -1751 2000
rect -1934 1848 -1871 1902
rect -1929 1847 -1871 1848
rect -1929 1838 -1907 1847
rect -1902 1838 -1871 1847
rect -1853 1894 -1847 1898
rect -1834 1896 -1799 1904
rect -1853 1890 -1841 1894
rect -1853 1884 -1837 1890
rect -1828 1886 -1824 1896
rect -1812 1886 -1808 1896
rect -1853 1873 -1834 1884
rect -1853 1867 -1828 1873
rect -1820 1872 -1816 1876
rect -1804 1873 -1800 1876
rect -1820 1868 -1811 1872
rect -1804 1868 -1801 1873
rect -1853 1856 -1834 1867
rect -1820 1864 -1816 1868
rect -1804 1864 -1800 1868
rect -1853 1850 -1837 1856
rect -1853 1846 -1841 1850
rect -1828 1849 -1824 1859
rect -1812 1849 -1808 1859
rect -1853 1842 -1847 1846
rect -1834 1841 -1799 1849
rect -1781 1739 -1751 1894
rect -1934 1683 -1871 1737
rect -1929 1682 -1871 1683
rect -1929 1673 -1907 1682
rect -1902 1673 -1871 1682
rect -1853 1729 -1847 1733
rect -1834 1731 -1799 1739
rect -1853 1725 -1841 1729
rect -1853 1719 -1837 1725
rect -1829 1721 -1825 1731
rect -1813 1721 -1809 1731
rect -1853 1708 -1836 1719
rect -1853 1702 -1829 1708
rect -1821 1707 -1817 1711
rect -1821 1703 -1812 1707
rect -1853 1691 -1836 1702
rect -1821 1699 -1817 1703
rect -1805 1699 -1801 1711
rect -1853 1685 -1837 1691
rect -1853 1681 -1841 1685
rect -1829 1684 -1825 1694
rect -1813 1684 -1809 1694
rect -1781 1689 -1751 1731
rect -1853 1677 -1847 1681
rect -1834 1676 -1799 1684
rect -1935 1448 -1872 1502
rect -1930 1447 -1872 1448
rect -1930 1438 -1908 1447
rect -1903 1438 -1872 1447
rect -1935 1191 -1872 1245
rect -1930 1190 -1872 1191
rect -1930 1181 -1908 1190
rect -1903 1181 -1872 1190
rect -1781 1199 -1751 1659
rect -1781 953 -1751 1169
rect -1935 897 -1872 951
rect -1930 896 -1872 897
rect -1930 887 -1908 896
rect -1903 887 -1872 896
rect -1854 943 -1848 947
rect -1835 945 -1800 953
rect -1854 939 -1842 943
rect -1854 933 -1838 939
rect -1829 935 -1825 945
rect -1813 935 -1809 945
rect -1854 922 -1835 933
rect -1854 916 -1829 922
rect -1821 921 -1817 925
rect -1821 917 -1812 921
rect -1854 905 -1835 916
rect -1821 913 -1817 917
rect -1805 913 -1801 925
rect -1854 899 -1838 905
rect -1854 895 -1842 899
rect -1829 898 -1825 908
rect -1813 898 -1809 908
rect -1854 891 -1848 895
rect -1835 890 -1800 898
rect -1781 719 -1751 945
rect -2403 651 -2339 705
rect -2398 650 -2339 651
rect -2398 641 -2376 650
rect -2371 641 -2339 650
rect -2323 695 -2321 697
rect -2323 687 -2302 695
rect -2323 649 -2321 687
rect -1781 650 -1751 689
rect -2403 335 -2339 389
rect -2398 334 -2339 335
rect -2398 325 -2376 334
rect -2371 325 -2339 334
rect -2323 357 -2304 365
rect -1815 359 -1812 364
rect -1781 334 -1751 642
rect -1781 249 -1751 326
rect -1781 -1 -1751 219
rect -1781 -181 -1751 -31
rect -1721 2319 -1631 2349
rect -1601 2319 -1391 2349
rect -1361 2319 -1151 2349
rect -1121 2319 -911 2349
rect -881 2319 -671 2349
rect -641 2319 -431 2349
rect -401 2319 -191 2349
rect -161 2319 258 2349
rect 288 2319 589 2349
rect 619 2319 849 2349
rect 879 2319 949 2349
rect -1721 2259 -1691 2319
rect -1721 1779 -1691 2229
rect -1721 1289 -1691 1749
rect -1721 809 -1691 1259
rect -1721 339 -1691 779
rect -1721 59 -1691 309
rect -1721 -121 -1691 29
rect -1661 2259 -1481 2289
rect -1451 2259 -1241 2289
rect -1211 2259 -1001 2289
rect -971 2259 -761 2289
rect -731 2259 -488 2289
rect -458 2259 -281 2289
rect -251 2259 178 2289
rect 208 2259 526 2289
rect 556 2259 759 2289
rect 789 2259 889 2289
rect -1661 1629 -1631 2259
rect 799 2229 829 2230
rect -1661 1139 -1631 1599
rect -1661 659 -1631 1109
rect -1661 189 -1631 629
rect -1661 -61 -1631 159
rect -1601 2199 -1331 2229
rect -1301 2199 -1091 2229
rect -1061 2199 -851 2229
rect -821 2199 -611 2229
rect -581 2199 -371 2229
rect -341 2199 107 2229
rect 137 2199 437 2229
rect 467 2199 669 2229
rect 699 2199 829 2229
rect -1601 1719 -1571 2169
rect -1601 1229 -1571 1689
rect -1601 749 -1571 1199
rect -1601 279 -1571 719
rect 799 2140 829 2199
rect 799 1972 829 2110
rect 799 1722 829 1942
rect 799 1472 829 1692
rect 799 1222 829 1442
rect 799 972 829 1192
rect 799 722 829 942
rect 243 558 249 596
rect -682 509 -677 516
rect -470 509 -468 516
rect -678 501 -677 509
rect -525 506 -510 508
rect -525 504 -500 506
rect -517 500 -500 504
rect -365 508 -364 517
rect -317 509 -313 513
rect -102 495 -74 500
rect -515 410 -500 414
rect -300 412 -230 418
rect -218 412 -216 418
rect -305 291 -242 297
rect -517 285 -499 291
rect -1601 -1 -1571 249
rect 799 513 829 692
rect 799 231 829 483
rect -1236 198 -1229 199
rect -1236 182 -1229 190
rect 799 -1 829 201
rect -1601 -31 -1569 -1
rect -1539 -31 -1329 -1
rect -1299 -31 -1089 -1
rect -1059 -31 -609 -1
rect -579 -31 -369 -1
rect -339 -31 89 -1
rect 119 -31 339 -1
rect 369 -31 671 -1
rect 701 -31 829 -1
rect 859 1881 889 2259
rect 859 1651 889 1851
rect 859 1381 889 1621
rect 859 1150 889 1351
rect 859 863 889 1120
rect 859 426 889 833
rect 859 199 889 396
rect -1257 -61 -1250 -59
rect -1180 -61 -1173 -58
rect -1029 -61 -1022 -59
rect -723 -61 -716 -59
rect 859 -61 889 169
rect -1631 -91 -1480 -61
rect -1450 -91 -1240 -61
rect -1210 -91 -1000 -61
rect -970 -91 -760 -61
rect -730 -91 -520 -61
rect -490 -91 -280 -61
rect -250 -91 -62 -61
rect -32 -91 188 -61
rect 218 -91 760 -61
rect 790 -91 889 -61
rect 919 2200 949 2319
rect 919 2032 949 2170
rect 919 1782 949 2002
rect 919 1532 949 1752
rect 919 1282 949 1502
rect 919 1032 949 1252
rect 919 782 949 1002
rect 919 573 949 752
rect 919 291 949 543
rect 919 101 949 261
rect -799 -93 -792 -91
rect 919 -121 949 71
rect -1721 -151 -1629 -121
rect -1599 -151 -1389 -121
rect -1359 -151 -1149 -121
rect -1119 -151 -909 -121
rect -879 -151 -669 -121
rect -639 -151 -429 -121
rect -399 -151 -189 -121
rect -159 -151 29 -121
rect 59 -151 279 -121
rect 309 -151 859 -121
rect 889 -151 949 -121
rect 979 2144 1009 2379
rect 979 1944 1009 2114
rect 979 1443 1009 1914
rect 1094 1790 1128 1799
rect 1133 1790 1155 1799
rect 1094 1789 1155 1790
rect 1094 1735 1160 1789
rect 979 1214 1009 1413
rect 979 680 1009 1184
rect 1093 1137 1128 1146
rect 1133 1137 1155 1146
rect 1093 1136 1155 1137
rect 1093 1082 1160 1136
rect 979 475 1009 650
rect 1034 643 1069 651
rect 1082 646 1088 650
rect 1043 633 1047 643
rect 1059 633 1063 643
rect 1076 642 1088 646
rect 1072 636 1088 642
rect 1035 627 1039 628
rect 1036 618 1039 627
rect 1051 624 1055 628
rect 1069 625 1088 636
rect 1046 620 1055 624
rect 1035 616 1039 618
rect 1051 616 1055 620
rect 1063 619 1088 625
rect 1069 608 1088 619
rect 1043 596 1047 606
rect 1059 596 1063 606
rect 1072 602 1088 608
rect 1076 598 1088 602
rect 1034 589 1069 596
rect 1082 594 1088 598
rect 1106 645 1137 654
rect 1142 645 1164 654
rect 1106 644 1164 645
rect 1106 590 1169 644
rect 979 376 1009 461
rect 1072 460 1082 470
rect 1599 388 1603 410
rect 1570 377 1603 388
rect 1599 362 1603 377
rect 1619 409 1651 418
rect 1656 409 1678 418
rect 1619 408 1678 409
rect 1619 354 1683 408
rect 979 214 1009 346
rect 1028 321 1038 332
rect 1050 321 1077 332
rect 979 31 1009 184
rect 1596 136 1600 156
rect 1059 125 1069 131
rect 1561 125 1600 136
rect 1595 124 1600 125
rect 1596 108 1600 124
rect 1616 155 1648 164
rect 1653 155 1675 164
rect 1616 154 1675 155
rect 1616 100 1680 154
rect 979 -181 1009 1
rect -1751 -211 -1540 -181
rect -1510 -211 -1379 -181
rect -1365 -211 -1300 -181
rect -1270 -211 -1160 -181
rect -1146 -211 -1060 -181
rect -1030 -211 -820 -181
rect -790 -211 -580 -181
rect -550 -211 -340 -181
rect -310 -211 -122 -181
rect -92 -211 128 -181
rect 158 -211 700 -181
rect 730 -211 1009 -181
rect -1316 -226 -1315 -219
rect -1324 -230 -1315 -226
rect -1114 -232 -1110 -216
rect -1119 -237 -1110 -232
rect 184 -250 191 -241
rect 211 -243 213 -242
rect 222 -243 223 -242
rect 211 -246 223 -243
rect 184 -254 201 -250
rect 238 -250 246 -241
rect 184 -266 191 -254
rect 215 -258 219 -253
rect 228 -254 246 -250
rect 211 -262 223 -258
rect -945 -297 -881 -266
rect -945 -302 -890 -297
rect -945 -324 -881 -302
rect -945 -329 -891 -324
rect -446 -297 -382 -266
rect 184 -270 201 -266
rect 238 -266 246 -254
rect 228 -270 246 -266
rect 184 -276 191 -270
rect 214 -276 220 -270
rect 238 -276 246 -270
rect 203 -279 231 -276
rect 197 -283 237 -279
rect 193 -289 241 -283
rect -446 -302 -391 -297
rect 189 -295 245 -289
rect -446 -324 -382 -302
rect -446 -329 -392 -324
rect 185 -344 249 -313
rect 185 -349 240 -344
rect 185 -371 249 -349
rect 185 -376 239 -371
rect -1409 -742 -1402 -720
rect -1202 -742 -1195 -724
rect -1423 -746 -1375 -742
rect -1219 -745 -1171 -742
rect -1431 -794 -1367 -762
rect -1431 -799 -1376 -794
rect -1431 -821 -1367 -799
rect -1431 -826 -1377 -821
rect -1227 -793 -1163 -761
rect -1227 -798 -1172 -793
rect -1227 -820 -1163 -798
rect -1227 -825 -1173 -820
<< metal2 >>
rect -1496 3041 -1442 3046
rect -1506 3040 -1442 3041
rect -1497 3035 -1442 3040
rect -1506 3019 -1442 3035
rect -1497 3014 -1442 3019
rect -1506 3013 -1442 3014
rect -1497 3008 -1442 3013
rect -1506 2982 -1442 3008
rect -1281 3041 -1227 3046
rect -1291 3040 -1227 3041
rect -1282 3035 -1227 3040
rect -1291 3019 -1227 3035
rect -1282 3014 -1227 3019
rect -1291 3013 -1227 3014
rect -1282 3008 -1227 3013
rect -1291 2982 -1227 3008
rect -1028 2567 -974 2572
rect -1038 2566 -974 2567
rect -1029 2561 -974 2566
rect -1038 2545 -974 2561
rect -1029 2540 -974 2545
rect -1038 2539 -974 2540
rect -1029 2534 -974 2539
rect -1038 2509 -974 2534
rect -781 2567 -727 2572
rect -791 2566 -727 2567
rect -782 2561 -727 2566
rect -791 2545 -727 2561
rect -782 2540 -727 2545
rect -791 2539 -727 2540
rect -782 2534 -727 2539
rect -791 2509 -727 2534
rect -563 2569 -509 2574
rect -573 2568 -509 2569
rect -564 2563 -509 2568
rect -573 2547 -509 2563
rect -564 2542 -509 2547
rect -573 2541 -509 2542
rect -564 2536 -509 2541
rect -573 2510 -509 2536
rect -289 2570 -235 2575
rect -299 2569 -235 2570
rect -290 2564 -235 2569
rect -299 2548 -235 2564
rect -290 2543 -235 2548
rect -299 2542 -235 2543
rect -290 2537 -235 2542
rect -299 2511 -235 2537
rect -1035 2426 -1027 2430
rect -788 2426 -780 2430
rect -1751 2379 -1661 2409
rect -1631 2379 -1527 2409
rect -1497 2379 -1421 2409
rect -1391 2379 -1301 2409
rect -1271 2379 -1181 2409
rect -1151 2379 -1061 2409
rect -1031 2379 -982 2409
rect -970 2379 -941 2409
rect -911 2379 -849 2409
rect -818 2379 -735 2409
rect -723 2379 -701 2409
rect -671 2379 -581 2409
rect -551 2379 -461 2409
rect -431 2379 -341 2409
rect -311 2379 -221 2409
rect -191 2379 0 2409
rect 30 2379 207 2409
rect 237 2379 321 2409
rect 351 2379 427 2409
rect 457 2379 699 2409
rect 729 2379 819 2409
rect 849 2379 939 2409
rect 969 2379 1009 2409
rect -1781 2289 -1751 2379
rect -2405 2052 -2341 2106
rect -2400 2051 -2341 2052
rect -2400 2042 -2399 2051
rect -2394 2042 -2378 2051
rect -2373 2042 -2372 2051
rect -2367 2042 -2341 2051
rect -1781 2015 -1751 2259
rect -1781 1906 -1751 2000
rect -1934 1848 -1871 1902
rect -1929 1847 -1871 1848
rect -1929 1838 -1928 1847
rect -1923 1838 -1907 1847
rect -1902 1838 -1901 1847
rect -1896 1838 -1871 1847
rect -1781 1809 -1751 1894
rect -1781 1739 -1751 1779
rect -1934 1683 -1871 1737
rect -1929 1682 -1871 1683
rect -1929 1673 -1928 1682
rect -1923 1673 -1907 1682
rect -1902 1673 -1901 1682
rect -1896 1673 -1871 1682
rect -1781 1689 -1751 1731
rect -1935 1448 -1872 1502
rect -1930 1447 -1872 1448
rect -1930 1438 -1929 1447
rect -1924 1438 -1908 1447
rect -1903 1438 -1902 1447
rect -1897 1438 -1872 1447
rect -1781 1319 -1751 1659
rect -1935 1191 -1872 1245
rect -1930 1190 -1872 1191
rect -1930 1181 -1929 1190
rect -1924 1181 -1908 1190
rect -1903 1181 -1902 1190
rect -1897 1181 -1872 1190
rect -1781 1199 -1751 1289
rect -1781 953 -1751 1169
rect -1935 897 -1872 951
rect -1930 896 -1872 897
rect -1930 887 -1929 896
rect -1924 887 -1908 896
rect -1903 887 -1902 896
rect -1897 887 -1872 896
rect -1781 839 -1751 945
rect -1781 719 -1751 809
rect -2403 651 -2339 705
rect -2398 650 -2339 651
rect -2398 641 -2397 650
rect -2392 641 -2376 650
rect -2371 641 -2370 650
rect -2365 641 -2339 650
rect -1781 650 -1751 689
rect -2403 335 -2339 389
rect -2398 334 -2339 335
rect -2398 325 -2397 334
rect -2392 325 -2376 334
rect -2371 325 -2370 334
rect -2365 325 -2339 334
rect -1781 369 -1751 642
rect -1781 334 -1751 339
rect -1781 249 -1751 326
rect -1781 89 -1751 219
rect -1781 -1 -1751 59
rect -1781 -75 -1751 -31
rect -1781 -181 -1751 -105
rect -1691 2319 -1631 2349
rect -1601 2319 -1511 2349
rect -1481 2319 -1391 2349
rect -1361 2319 -1297 2349
rect -1267 2319 -1151 2349
rect -1121 2319 -911 2349
rect -881 2319 -848 2349
rect -818 2319 -671 2349
rect -641 2319 -551 2349
rect -521 2319 -431 2349
rect -401 2319 -311 2349
rect -281 2319 -191 2349
rect -161 2319 -62 2349
rect -32 2319 138 2349
rect 168 2319 258 2349
rect 288 2319 431 2349
rect 461 2319 589 2349
rect 619 2319 729 2349
rect 759 2319 849 2349
rect 879 2319 949 2349
rect -1721 2259 -1691 2319
rect -1721 1779 -1691 2229
rect -1721 1659 -1691 1749
rect -1721 1289 -1691 1629
rect -1721 1169 -1691 1259
rect -1721 809 -1691 1139
rect -1721 689 -1691 779
rect -1721 339 -1691 659
rect -1721 219 -1691 309
rect -1721 59 -1691 189
rect -1721 -33 -1691 29
rect -1721 -121 -1691 -63
rect -1661 2259 -1601 2289
rect -1571 2259 -1481 2289
rect -1451 2259 -1361 2289
rect -1331 2259 -1241 2289
rect -1211 2259 -1121 2289
rect -1091 2259 -1001 2289
rect -971 2259 -881 2289
rect -851 2259 -761 2289
rect -731 2259 -641 2289
rect -611 2259 -488 2289
rect -458 2259 -401 2289
rect -371 2259 -281 2289
rect -251 2259 -132 2289
rect -102 2259 54 2289
rect 84 2259 178 2289
rect 208 2259 377 2289
rect 407 2259 526 2289
rect 556 2259 642 2289
rect 669 2259 759 2289
rect 789 2259 889 2289
rect -1661 2229 -1631 2259
rect 799 2229 829 2230
rect -1661 1749 -1631 2199
rect -1661 1629 -1631 1719
rect -1661 1294 -1631 1599
rect -1661 1139 -1631 1264
rect -1661 779 -1631 1109
rect -1661 659 -1631 749
rect -1661 309 -1631 629
rect -1661 189 -1631 279
rect -1661 29 -1631 159
rect -1661 -61 -1631 -1
rect -1601 2199 -1451 2229
rect -1421 2199 -1331 2229
rect -1301 2199 -1211 2229
rect -1181 2199 -1091 2229
rect -1061 2199 -971 2229
rect -941 2199 -851 2229
rect -821 2199 -731 2229
rect -701 2199 -611 2229
rect -581 2199 -491 2229
rect -461 2199 -371 2229
rect -341 2199 -221 2229
rect -191 2199 -6 2229
rect 24 2199 107 2229
rect 137 2199 259 2229
rect 289 2199 437 2229
rect 467 2199 559 2229
rect 589 2199 669 2229
rect 699 2199 789 2229
rect 819 2199 829 2229
rect -1601 1719 -1571 2169
rect -1601 1599 -1571 1689
rect -1601 1229 -1571 1569
rect -1601 1109 -1571 1199
rect -1601 749 -1571 1079
rect -1601 629 -1571 719
rect 799 2140 829 2199
rect 799 2069 829 2110
rect 799 1972 829 2039
rect 799 1910 829 1942
rect 799 1722 829 1880
rect 799 1611 829 1692
rect 799 1472 829 1581
rect 799 1344 829 1442
rect 799 1222 829 1314
rect 799 1115 829 1192
rect 799 972 829 1085
rect 799 722 829 942
rect 799 631 829 692
rect -1601 279 -1571 599
rect 799 513 829 601
rect -1601 159 -1571 249
rect 218 240 219 252
rect 799 231 829 483
rect -1601 -1 -1571 129
rect 799 -1 829 201
rect -1601 -31 -1569 -1
rect -1539 -31 -1450 -1
rect -1420 -31 -1329 -1
rect -1299 -31 -1210 -1
rect -1180 -31 -1089 -1
rect -1059 -31 -970 -1
rect -940 -31 -730 -1
rect -700 -31 -609 -1
rect -579 -31 -490 -1
rect -460 -31 -369 -1
rect -339 -31 -250 -1
rect -220 -31 -32 -1
rect -2 -31 89 -1
rect 119 -31 218 -1
rect 248 -31 339 -1
rect 369 -31 671 -1
rect 701 -31 790 -1
rect 820 -31 829 -1
rect 859 2170 889 2259
rect 859 2002 889 2140
rect 859 1881 889 1972
rect 859 1752 889 1851
rect 859 1651 889 1722
rect 859 1502 889 1621
rect 859 1381 889 1472
rect 859 1252 889 1351
rect 859 1150 889 1222
rect 859 1002 889 1120
rect 859 863 889 972
rect 859 752 889 833
rect 859 543 889 722
rect 859 426 889 513
rect 859 261 889 396
rect 859 199 889 231
rect 859 71 889 169
rect -1257 -61 -1250 -59
rect -1180 -61 -1173 -58
rect -1029 -61 -1022 -59
rect -723 -61 -716 -59
rect 859 -61 889 41
rect -1631 -91 -1599 -61
rect -1569 -91 -1480 -61
rect -1450 -91 -1359 -61
rect -1329 -91 -1240 -61
rect -1210 -91 -1119 -61
rect -1089 -91 -1000 -61
rect -970 -91 -879 -61
rect -849 -91 -760 -61
rect -730 -91 -639 -61
rect -609 -91 -520 -61
rect -490 -91 -280 -61
rect -250 -91 -62 -61
rect -32 -91 59 -61
rect 89 -91 188 -61
rect 218 -91 309 -61
rect 339 -91 642 -61
rect 671 -91 760 -61
rect 790 -91 889 -61
rect 919 2200 949 2319
rect 919 2148 949 2170
rect 919 2032 949 2118
rect 919 1782 949 2002
rect 919 1685 949 1752
rect 919 1532 949 1655
rect 919 1414 949 1502
rect 919 1282 949 1384
rect 919 1182 949 1252
rect 919 1032 949 1152
rect 919 782 949 1002
rect 919 624 949 752
rect 919 573 949 594
rect 919 467 949 543
rect 919 291 949 437
rect 919 101 949 261
rect 919 -32 949 71
rect -799 -93 -792 -91
rect 919 -121 949 -62
rect -1721 -151 -1629 -121
rect -1599 -151 -1510 -121
rect -1480 -151 -1389 -121
rect -1359 -151 -1270 -121
rect -1240 -151 -1149 -121
rect -1119 -151 -1030 -121
rect -1000 -151 -909 -121
rect -879 -151 -790 -121
rect -760 -151 -669 -121
rect -639 -151 -550 -121
rect -520 -151 -429 -121
rect -399 -151 -310 -121
rect -280 -151 -189 -121
rect -159 -151 -92 -121
rect -62 -151 29 -121
rect 59 -151 158 -121
rect 188 -151 279 -121
rect 309 -151 730 -121
rect 760 -151 859 -121
rect 889 -151 949 -121
rect 979 2230 1009 2379
rect 979 2144 1009 2200
rect 979 2062 1009 2114
rect 979 1944 1009 2032
rect 979 1812 1009 1914
rect 979 1562 1009 1782
rect 1094 1790 1122 1799
rect 1127 1790 1128 1799
rect 1133 1790 1149 1799
rect 1154 1790 1155 1799
rect 1094 1789 1155 1790
rect 1094 1735 1160 1789
rect 979 1443 1009 1532
rect 979 1312 1009 1413
rect 979 1214 1009 1282
rect 979 1062 1009 1184
rect 1093 1137 1122 1146
rect 1127 1137 1128 1146
rect 1133 1137 1149 1146
rect 1154 1137 1155 1146
rect 1093 1136 1155 1137
rect 1093 1082 1160 1136
rect 979 812 1009 1032
rect 979 680 1009 782
rect 979 603 1009 650
rect 1106 645 1131 654
rect 1136 645 1137 654
rect 1142 645 1158 654
rect 1163 645 1164 654
rect 1106 644 1164 645
rect 1106 590 1169 644
rect 979 475 1009 573
rect 979 376 1009 461
rect 1619 409 1645 418
rect 1650 409 1651 418
rect 1656 409 1672 418
rect 1677 409 1678 418
rect 1619 408 1678 409
rect 1619 354 1683 408
rect 979 321 1009 346
rect 979 214 1009 291
rect 979 131 1009 184
rect 1616 155 1642 164
rect 1647 155 1648 164
rect 1653 155 1669 164
rect 1674 155 1675 164
rect 1616 154 1675 155
rect 979 31 1009 101
rect 1616 100 1680 154
rect 979 -181 1009 1
rect -1751 -211 -1660 -181
rect -1630 -211 -1540 -181
rect -1510 -211 -1420 -181
rect -1390 -211 -1379 -181
rect -1365 -211 -1300 -181
rect -1270 -211 -1207 -181
rect -1177 -211 -1160 -181
rect -1146 -211 -1060 -181
rect -1030 -211 -940 -181
rect -910 -211 -820 -181
rect -790 -211 -700 -181
rect -670 -211 -580 -181
rect -550 -211 -460 -181
rect -430 -211 -340 -181
rect -310 -211 -220 -181
rect -190 -211 -122 -181
rect -92 -211 -2 -181
rect 28 -211 128 -181
rect 158 -211 248 -181
rect 278 -211 700 -181
rect 730 -211 918 -181
rect 948 -211 1009 -181
rect -945 -291 -881 -266
rect -945 -296 -890 -291
rect -945 -297 -881 -296
rect -945 -302 -890 -297
rect -945 -318 -881 -302
rect -945 -323 -890 -318
rect -945 -324 -881 -323
rect -945 -329 -891 -324
rect -446 -291 -382 -266
rect -446 -296 -391 -291
rect -446 -297 -382 -296
rect -446 -302 -391 -297
rect -446 -318 -382 -302
rect -446 -323 -391 -318
rect -446 -324 -382 -323
rect -446 -329 -392 -324
rect 185 -338 249 -313
rect 185 -343 240 -338
rect 185 -344 249 -343
rect 185 -349 240 -344
rect 185 -365 249 -349
rect 185 -370 240 -365
rect 185 -371 249 -370
rect 185 -376 239 -371
rect -1431 -788 -1367 -762
rect -1431 -793 -1376 -788
rect -1431 -794 -1367 -793
rect -1431 -799 -1376 -794
rect -1431 -815 -1367 -799
rect -1431 -820 -1376 -815
rect -1431 -821 -1367 -820
rect -1431 -826 -1377 -821
rect -1227 -787 -1163 -761
rect -1227 -792 -1172 -787
rect -1227 -793 -1163 -792
rect -1227 -798 -1172 -793
rect -1227 -814 -1163 -798
rect -1227 -819 -1172 -814
rect -1227 -820 -1163 -819
rect -1227 -825 -1173 -820
<< m123contact >>
rect -1506 3041 -1496 3046
rect -1506 3014 -1497 3019
rect -1291 3041 -1281 3046
rect -1291 3014 -1282 3019
rect -1504 2966 -1444 2972
rect -1289 2966 -1229 2972
rect -1038 2567 -1028 2572
rect -1038 2540 -1029 2545
rect -791 2567 -781 2572
rect -791 2540 -782 2545
rect -573 2569 -563 2574
rect -573 2542 -564 2547
rect -299 2570 -289 2575
rect -299 2543 -290 2548
rect -1034 2491 -978 2497
rect -787 2491 -731 2497
rect -1558 2441 -1547 2452
rect -1486 2438 -1463 2449
rect -1418 2429 -1408 2442
rect -1340 2439 -1331 2450
rect -1253 2432 -1243 2445
rect -1201 2434 -1191 2448
rect -1035 2430 -1027 2437
rect -1008 2432 -1003 2439
rect -980 2432 -972 2437
rect -788 2430 -780 2437
rect -761 2433 -756 2438
rect -733 2432 -725 2437
rect -1781 2379 -1751 2409
rect -1527 2379 -1497 2409
rect -1301 2379 -1271 2409
rect -1061 2379 -1031 2409
rect -982 2379 -970 2414
rect -849 2379 -818 2409
rect -735 2379 -723 2409
rect -581 2379 -551 2409
rect -341 2379 -311 2409
rect 321 2379 351 2409
rect 699 2379 729 2409
rect 939 2379 969 2409
rect -1814 2135 -1801 2147
rect -2405 2042 -2400 2052
rect -2378 2042 -2373 2051
rect -2331 2044 -2325 2104
rect -1816 2082 -1808 2093
rect -1815 1997 -1807 2005
rect -1781 2000 -1751 2015
rect -1934 1838 -1929 1848
rect -1907 1838 -1902 1847
rect -1859 1842 -1853 1898
rect -1799 1896 -1791 1904
rect -1781 1894 -1751 1906
rect -1801 1868 -1796 1873
rect -1799 1841 -1793 1849
rect -1934 1673 -1929 1683
rect -1907 1673 -1902 1682
rect -1859 1677 -1853 1733
rect -1799 1731 -1791 1739
rect -1781 1731 -1751 1739
rect -1801 1703 -1796 1708
rect -1799 1676 -1793 1684
rect -1781 1659 -1751 1689
rect -1935 1438 -1930 1448
rect -1908 1438 -1903 1447
rect -1935 1181 -1930 1191
rect -1908 1181 -1903 1190
rect -1781 1169 -1751 1199
rect -1935 887 -1930 897
rect -1908 887 -1903 896
rect -1860 891 -1854 947
rect -1800 945 -1792 953
rect -1781 945 -1751 953
rect -1801 917 -1795 923
rect -1800 890 -1794 898
rect -1808 742 -1800 750
rect -2403 641 -2398 651
rect -2376 641 -2371 650
rect -2329 643 -2323 703
rect -1806 690 -1800 696
rect -1781 689 -1751 719
rect -1781 642 -1751 650
rect -1807 604 -1800 612
rect -1809 411 -1797 418
rect -2403 325 -2398 335
rect -2376 325 -2371 334
rect -2329 327 -2323 387
rect -1812 359 -1804 364
rect -1781 326 -1751 334
rect -1813 272 -1797 280
rect -1781 219 -1751 249
rect -1781 -31 -1751 -1
rect -1631 2319 -1601 2349
rect -1391 2319 -1361 2349
rect -1151 2319 -1121 2349
rect -911 2319 -881 2349
rect -671 2319 -641 2349
rect -431 2319 -401 2349
rect -191 2319 -161 2349
rect 258 2319 288 2349
rect 589 2319 619 2349
rect 849 2319 879 2349
rect -1721 2229 -1691 2259
rect -1721 1749 -1691 1779
rect -1721 1259 -1691 1289
rect -1721 779 -1691 809
rect -1721 309 -1691 339
rect -1721 29 -1691 59
rect -1481 2259 -1451 2289
rect -1241 2259 -1211 2289
rect -1001 2259 -971 2289
rect -761 2259 -731 2289
rect -488 2259 -458 2289
rect -281 2259 -251 2289
rect 178 2259 208 2289
rect 526 2259 556 2289
rect 759 2259 789 2289
rect -1661 1599 -1631 1629
rect -1661 1109 -1631 1139
rect -1661 629 -1631 659
rect -1661 159 -1631 189
rect -1331 2199 -1301 2229
rect -1091 2199 -1061 2229
rect -851 2199 -821 2229
rect -611 2199 -581 2229
rect -371 2199 -341 2229
rect 107 2199 137 2229
rect 437 2199 467 2229
rect 669 2199 699 2229
rect -1601 2169 -1571 2199
rect -1601 1689 -1571 1719
rect -1601 1199 -1571 1229
rect -1601 719 -1571 749
rect 799 2110 829 2140
rect 799 1942 829 1972
rect 799 1692 829 1722
rect 799 1442 829 1472
rect 799 1192 829 1222
rect 799 942 829 972
rect 799 692 829 722
rect 242 596 249 605
rect -285 550 -278 556
rect -686 501 -678 509
rect -632 501 -625 509
rect -582 503 -572 509
rect -500 500 -494 506
rect -472 501 -464 509
rect -420 501 -412 509
rect -367 499 -358 508
rect -321 501 -312 509
rect -74 495 -67 502
rect 799 483 829 513
rect -500 410 -495 415
rect -230 412 -218 424
rect -499 285 -491 291
rect -242 288 -230 300
rect -1601 249 -1571 279
rect 213 240 218 252
rect 243 202 248 209
rect 265 208 275 218
rect 799 201 829 231
rect -1314 190 -1305 198
rect -1238 190 -1229 198
rect -1255 181 -1248 187
rect -1177 180 -1170 186
rect -1161 184 -1153 192
rect -1085 183 -1077 191
rect -1027 181 -1020 187
rect -1010 183 -1002 191
rect -950 182 -943 188
rect -934 181 -926 189
rect -857 185 -849 193
rect -798 180 -791 186
rect -780 184 -772 192
rect -721 179 -713 186
rect -522 168 -514 174
rect -1569 -31 -1539 -1
rect -1329 -31 -1299 -1
rect -1089 -31 -1059 -1
rect -609 -31 -579 -1
rect -369 -31 -339 -1
rect 89 -31 119 -1
rect 339 -31 369 -1
rect 671 -31 701 -1
rect 859 1851 889 1881
rect 859 1621 889 1651
rect 859 1351 889 1381
rect 859 1120 889 1150
rect 859 833 889 863
rect 859 396 889 426
rect 859 169 889 199
rect -1661 -91 -1631 -61
rect -1480 -91 -1450 -61
rect -1240 -91 -1210 -61
rect -1000 -91 -970 -61
rect -760 -91 -730 -61
rect -520 -91 -490 -61
rect -280 -91 -250 -61
rect -62 -91 -32 -61
rect 188 -91 218 -61
rect 760 -91 790 -61
rect 919 2170 949 2200
rect 919 2002 949 2032
rect 919 1752 949 1782
rect 919 1502 949 1532
rect 919 1252 949 1282
rect 919 1002 949 1032
rect 919 752 949 782
rect 919 543 949 573
rect 919 261 949 291
rect 919 71 949 101
rect -1629 -151 -1599 -121
rect -1389 -151 -1359 -121
rect -1149 -151 -1119 -121
rect -909 -151 -879 -121
rect -669 -151 -639 -121
rect -429 -151 -399 -121
rect -189 -151 -159 -121
rect 29 -151 59 -121
rect 279 -151 309 -121
rect 859 -151 889 -121
rect 979 2114 1009 2144
rect 979 1914 1009 1944
rect 1128 1790 1133 1799
rect 1155 1789 1160 1799
rect 979 1413 1009 1443
rect 979 1184 1009 1214
rect 1128 1137 1133 1146
rect 1155 1136 1160 1146
rect 979 650 1009 680
rect 1026 643 1034 651
rect 1027 618 1036 627
rect 1025 589 1034 596
rect 1088 594 1094 650
rect 1137 645 1142 654
rect 1164 644 1169 654
rect 979 461 1009 475
rect 1056 460 1072 476
rect 1069 376 1076 383
rect 979 346 1009 376
rect 1603 356 1609 416
rect 1651 409 1656 418
rect 1678 408 1683 418
rect 1038 321 1050 333
rect 979 184 1027 214
rect 1059 211 1068 218
rect 1051 125 1059 131
rect 1600 102 1606 162
rect 1648 155 1653 164
rect 1675 154 1680 164
rect 1057 73 1066 80
rect 979 1 1009 31
rect -1781 -211 -1751 -181
rect -1540 -211 -1510 -181
rect -1379 -211 -1365 -181
rect -1300 -211 -1270 -181
rect -1160 -211 -1146 -181
rect -1060 -211 -1030 -181
rect -820 -211 -790 -181
rect -580 -211 -550 -181
rect -340 -211 -310 -181
rect -122 -211 -92 -181
rect 128 -211 158 -181
rect 700 -211 730 -181
rect -1462 -229 -1454 -220
rect -1409 -231 -1400 -224
rect -1326 -226 -1316 -216
rect -1258 -227 -1248 -219
rect -1205 -232 -1198 -226
rect -1124 -232 -1114 -216
rect 184 -241 191 -232
rect 213 -243 222 -234
rect 238 -241 246 -233
rect -890 -302 -881 -297
rect -891 -329 -881 -324
rect -391 -302 -382 -297
rect 189 -301 245 -295
rect -392 -329 -382 -324
rect 240 -349 249 -344
rect 239 -376 249 -371
rect -1429 -752 -1369 -746
rect -1225 -751 -1165 -745
rect -1376 -799 -1367 -794
rect -1377 -826 -1367 -821
rect -1172 -798 -1163 -793
rect -1173 -825 -1163 -820
<< metal3 >>
rect -1496 3041 -1442 3046
rect -1506 3040 -1442 3041
rect -1497 3035 -1442 3040
rect -1506 3034 -1442 3035
rect -1497 3029 -1442 3034
rect -1506 3019 -1442 3029
rect -1497 3014 -1442 3019
rect -1506 3013 -1442 3014
rect -1497 3008 -1442 3013
rect -1506 3007 -1442 3008
rect -1497 3002 -1442 3007
rect -1506 2982 -1442 3002
rect -1281 3041 -1227 3046
rect -1291 3040 -1227 3041
rect -1282 3035 -1227 3040
rect -1291 3034 -1227 3035
rect -1282 3029 -1227 3034
rect -1291 3019 -1227 3029
rect -1282 3014 -1227 3019
rect -1291 3013 -1227 3014
rect -1282 3008 -1227 3013
rect -1291 3007 -1227 3008
rect -1282 3002 -1227 3007
rect -1291 2982 -1227 3002
rect -1028 2567 -974 2572
rect -1038 2566 -974 2567
rect -1029 2561 -974 2566
rect -1038 2560 -974 2561
rect -1029 2555 -974 2560
rect -1038 2545 -974 2555
rect -1029 2540 -974 2545
rect -1038 2539 -974 2540
rect -1029 2534 -974 2539
rect -1038 2533 -974 2534
rect -1029 2528 -974 2533
rect -1038 2509 -974 2528
rect -781 2567 -727 2572
rect -791 2566 -727 2567
rect -782 2561 -727 2566
rect -791 2560 -727 2561
rect -782 2555 -727 2560
rect -791 2545 -727 2555
rect -782 2540 -727 2545
rect -791 2539 -727 2540
rect -782 2534 -727 2539
rect -791 2533 -727 2534
rect -782 2528 -727 2533
rect -791 2509 -727 2528
rect -563 2569 -509 2574
rect -573 2568 -509 2569
rect -564 2563 -509 2568
rect -573 2562 -509 2563
rect -564 2557 -509 2562
rect -573 2547 -509 2557
rect -564 2542 -509 2547
rect -573 2541 -509 2542
rect -564 2536 -509 2541
rect -573 2535 -509 2536
rect -564 2530 -509 2535
rect -573 2510 -509 2530
rect -289 2570 -235 2575
rect -299 2569 -235 2570
rect -290 2564 -235 2569
rect -299 2563 -235 2564
rect -290 2558 -235 2563
rect -299 2548 -235 2558
rect -290 2543 -235 2548
rect -299 2542 -235 2543
rect -290 2537 -235 2542
rect -299 2536 -235 2537
rect -290 2531 -235 2536
rect -299 2511 -235 2531
rect -1558 2452 -1547 2454
rect -1340 2450 -1331 2451
rect -1558 2424 -1547 2441
rect -1560 2409 -1497 2424
rect -1340 2426 -1331 2439
rect -1341 2414 -1273 2426
rect -1341 2413 -1271 2414
rect -980 2427 -972 2432
rect -982 2414 -970 2427
rect -733 2427 -725 2432
rect -1301 2409 -1271 2413
rect -1751 2379 -1661 2409
rect -1631 2379 -1527 2409
rect -1497 2379 -1421 2409
rect -1391 2379 -1301 2409
rect -1271 2379 -1181 2409
rect -1151 2379 -1061 2409
rect -1031 2379 -982 2409
rect -735 2409 -723 2427
rect -970 2379 -941 2409
rect -911 2379 -849 2409
rect -818 2379 -735 2409
rect -723 2379 -701 2409
rect -671 2379 -581 2409
rect -551 2379 -461 2409
rect -431 2379 -341 2409
rect -311 2379 -221 2409
rect -191 2379 0 2409
rect 30 2379 207 2409
rect 237 2379 321 2409
rect 351 2379 427 2409
rect 457 2379 699 2409
rect 729 2379 819 2409
rect 849 2379 939 2409
rect 969 2379 1009 2409
rect -1781 2289 -1751 2379
rect -2405 2052 -2341 2106
rect -2400 2051 -2341 2052
rect -2400 2042 -2399 2051
rect -2394 2042 -2393 2051
rect -2388 2042 -2378 2051
rect -2373 2042 -2372 2051
rect -2367 2042 -2366 2051
rect -2361 2042 -2341 2051
rect -1781 2015 -1751 2259
rect -1807 2000 -1781 2015
rect -1807 1997 -1790 2000
rect -1781 1906 -1751 2000
rect -1934 1848 -1871 1902
rect -1929 1847 -1871 1848
rect -1929 1838 -1928 1847
rect -1923 1838 -1922 1847
rect -1917 1838 -1907 1847
rect -1902 1838 -1901 1847
rect -1896 1838 -1895 1847
rect -1890 1838 -1871 1847
rect -1791 1896 -1781 1904
rect -1781 1809 -1751 1894
rect -1781 1739 -1751 1779
rect -1934 1683 -1871 1737
rect -1929 1682 -1871 1683
rect -1929 1673 -1928 1682
rect -1923 1673 -1922 1682
rect -1917 1673 -1907 1682
rect -1902 1673 -1901 1682
rect -1896 1673 -1895 1682
rect -1890 1673 -1871 1682
rect -1791 1731 -1781 1739
rect -1781 1689 -1751 1731
rect -1935 1448 -1872 1502
rect -1930 1447 -1872 1448
rect -1930 1438 -1929 1447
rect -1924 1438 -1923 1447
rect -1918 1438 -1908 1447
rect -1903 1438 -1902 1447
rect -1897 1438 -1896 1447
rect -1891 1438 -1872 1447
rect -1781 1319 -1751 1659
rect -1935 1191 -1872 1245
rect -1930 1190 -1872 1191
rect -1930 1181 -1929 1190
rect -1924 1181 -1923 1190
rect -1918 1181 -1908 1190
rect -1903 1181 -1902 1190
rect -1897 1181 -1896 1190
rect -1891 1181 -1872 1190
rect -1781 1199 -1751 1289
rect -1781 953 -1751 1169
rect -1935 897 -1872 951
rect -1930 896 -1872 897
rect -1930 887 -1929 896
rect -1924 887 -1923 896
rect -1918 887 -1908 896
rect -1903 887 -1902 896
rect -1897 887 -1896 896
rect -1891 887 -1872 896
rect -1792 945 -1781 953
rect -1781 839 -1751 945
rect -1781 719 -1751 809
rect -2403 651 -2339 705
rect -2398 650 -2339 651
rect -2398 641 -2397 650
rect -2392 641 -2391 650
rect -2386 641 -2376 650
rect -2371 641 -2370 650
rect -2365 641 -2364 650
rect -2359 641 -2339 650
rect -1781 650 -1751 689
rect -1800 642 -1781 650
rect -1800 604 -1790 642
rect -2403 335 -2339 389
rect -2398 334 -2339 335
rect -2398 325 -2397 334
rect -2392 325 -2391 334
rect -2386 325 -2376 334
rect -2371 325 -2370 334
rect -2365 325 -2364 334
rect -2359 325 -2339 334
rect -1781 369 -1751 642
rect -1781 334 -1751 339
rect -1798 326 -1781 334
rect -1798 280 -1789 326
rect -1797 272 -1789 280
rect -1781 249 -1751 326
rect -1781 89 -1751 219
rect -1781 -1 -1751 59
rect -1781 -75 -1751 -31
rect -1781 -181 -1751 -105
rect -1691 2319 -1631 2349
rect -1601 2319 -1511 2349
rect -1481 2319 -1453 2349
rect -1439 2319 -1391 2349
rect -1361 2319 -1297 2349
rect -1267 2319 -1246 2349
rect -1216 2319 -1151 2349
rect -1121 2319 -1039 2349
rect -1023 2319 -911 2349
rect -881 2319 -848 2349
rect -818 2319 -792 2349
rect -776 2319 -671 2349
rect -641 2319 -551 2349
rect -521 2319 -431 2349
rect -401 2319 -311 2349
rect -281 2319 -191 2349
rect -161 2319 -62 2349
rect -32 2319 138 2349
rect 168 2319 258 2349
rect 288 2319 431 2349
rect 461 2319 589 2349
rect 619 2319 729 2349
rect 759 2319 849 2349
rect 879 2319 949 2349
rect -1721 2259 -1691 2319
rect -1721 2068 -1691 2229
rect -1721 1851 -1691 2055
rect -1721 1779 -1691 1839
rect -1721 1686 -1691 1749
rect -1721 1659 -1691 1674
rect -1721 1289 -1691 1629
rect -1721 1169 -1691 1259
rect -1721 900 -1691 1139
rect -1721 809 -1691 888
rect -1721 705 -1691 779
rect -1721 689 -1691 697
rect -1721 389 -1691 659
rect -1721 339 -1691 381
rect -1721 219 -1691 309
rect -1721 59 -1691 189
rect -1721 -33 -1691 29
rect -1721 -121 -1691 -63
rect -1661 2259 -1601 2289
rect -1571 2259 -1481 2289
rect -1451 2259 -1361 2289
rect -1331 2259 -1241 2289
rect -1211 2259 -1121 2289
rect -1091 2259 -1001 2289
rect -971 2259 -881 2289
rect -851 2259 -761 2289
rect -731 2259 -641 2289
rect -611 2259 -557 2289
rect -527 2259 -488 2289
rect -458 2259 -401 2289
rect -371 2259 -281 2289
rect -251 2259 -132 2289
rect -102 2259 54 2289
rect 84 2259 178 2289
rect 208 2259 377 2289
rect 407 2259 526 2289
rect 556 2259 642 2289
rect 669 2259 759 2289
rect 789 2259 889 2289
rect -1661 2229 -1631 2259
rect 799 2229 829 2230
rect -1661 1749 -1631 2199
rect -1661 1629 -1631 1719
rect -1661 1294 -1631 1599
rect -1661 1228 -1631 1264
rect -1661 1139 -1631 1198
rect -1661 779 -1631 1109
rect -1661 659 -1631 749
rect -1661 309 -1631 629
rect -1661 189 -1631 279
rect -1661 29 -1631 159
rect -1661 -61 -1631 -1
rect -1601 2199 -1451 2229
rect -1421 2199 -1331 2229
rect -1301 2199 -1211 2229
rect -1181 2199 -1091 2229
rect -1061 2199 -971 2229
rect -941 2199 -851 2229
rect -821 2199 -731 2229
rect -701 2199 -611 2229
rect -581 2199 -491 2229
rect -461 2199 -371 2229
rect -341 2199 -282 2229
rect -252 2199 -221 2229
rect -191 2199 -6 2229
rect 24 2199 107 2229
rect 137 2199 259 2229
rect 289 2199 437 2229
rect 467 2199 559 2229
rect 589 2199 669 2229
rect 699 2199 789 2229
rect 819 2199 829 2229
rect -1601 1719 -1571 2169
rect -1601 1599 -1571 1689
rect -1601 1485 -1571 1569
rect -1601 1229 -1571 1455
rect -1601 1109 -1571 1199
rect -1601 749 -1571 1079
rect -1601 629 -1571 719
rect 799 2140 829 2199
rect 799 2069 829 2110
rect 799 1972 829 2039
rect 799 1910 829 1942
rect 799 1722 829 1880
rect 799 1611 829 1692
rect 799 1472 829 1581
rect 799 1344 829 1442
rect 799 1222 829 1314
rect 799 1115 829 1192
rect 799 972 829 1085
rect 799 722 829 942
rect 799 631 829 692
rect -1601 279 -1571 599
rect 799 513 829 601
rect -1601 159 -1571 249
rect 218 240 219 252
rect 799 231 829 483
rect -1601 -1 -1571 129
rect 799 -1 829 201
rect -1601 -31 -1569 -1
rect -1539 -31 -1450 -1
rect -1420 -31 -1329 -1
rect -1299 -31 -1210 -1
rect -1180 -31 -1089 -1
rect -1059 -31 -970 -1
rect -940 -31 -928 -1
rect -898 -31 -730 -1
rect -700 -31 -609 -1
rect -579 -31 -490 -1
rect -460 -31 -369 -1
rect -339 -31 -250 -1
rect -220 -31 -32 -1
rect -2 -31 89 -1
rect 119 -31 218 -1
rect 248 -31 339 -1
rect 369 -31 671 -1
rect 701 -31 790 -1
rect 820 -31 829 -1
rect 859 2170 889 2259
rect 859 2002 889 2140
rect 859 1881 889 1972
rect 859 1752 889 1851
rect 859 1651 889 1722
rect 859 1502 889 1621
rect 859 1381 889 1472
rect 859 1252 889 1351
rect 859 1150 889 1222
rect 859 1002 889 1120
rect 859 863 889 972
rect 859 752 889 833
rect 859 543 889 722
rect 859 426 889 513
rect 859 261 889 396
rect 859 199 889 231
rect 859 71 889 169
rect -1257 -61 -1250 -59
rect -1180 -61 -1173 -58
rect -1029 -61 -1022 -59
rect -723 -61 -716 -59
rect 859 -61 889 41
rect -1631 -91 -1599 -61
rect -1569 -91 -1480 -61
rect -1450 -91 -1359 -61
rect -1329 -91 -1240 -61
rect -1210 -91 -1119 -61
rect -1089 -91 -1000 -61
rect -970 -91 -879 -61
rect -849 -91 -760 -61
rect -730 -91 -639 -61
rect -609 -91 -520 -61
rect -490 -91 -429 -61
rect -399 -91 -280 -61
rect -250 -91 -62 -61
rect -32 -91 59 -61
rect 89 -91 188 -61
rect 218 -91 309 -61
rect 339 -91 642 -61
rect 671 -91 760 -61
rect 790 -91 889 -61
rect 919 2200 949 2319
rect 919 2148 949 2170
rect 919 2080 949 2118
rect 919 2032 949 2067
rect 919 1782 949 2002
rect 919 1685 949 1752
rect 919 1532 949 1655
rect 919 1414 949 1502
rect 919 1282 949 1384
rect 919 1182 949 1252
rect 919 1130 949 1152
rect 919 1032 949 1100
rect 919 782 949 1002
rect 919 662 949 752
rect 919 624 949 632
rect 919 573 949 594
rect 919 467 949 543
rect 919 420 949 437
rect 919 291 949 407
rect 919 151 949 261
rect 919 101 949 138
rect 919 -32 949 71
rect -799 -93 -792 -91
rect 919 -121 949 -62
rect -1721 -151 -1629 -121
rect -1599 -151 -1510 -121
rect -1480 -151 -1433 -121
rect -1420 -151 -1389 -121
rect -1359 -151 -1270 -121
rect -1240 -151 -1214 -121
rect -1201 -151 -1149 -121
rect -1119 -151 -1030 -121
rect -1000 -151 -909 -121
rect -879 -151 -790 -121
rect -760 -151 -669 -121
rect -639 -151 -550 -121
rect -520 -151 -429 -121
rect -399 -151 -310 -121
rect -280 -151 -189 -121
rect -159 -151 -92 -121
rect -62 -151 29 -121
rect 59 -151 158 -121
rect 188 -151 279 -121
rect 309 -151 730 -121
rect 760 -151 859 -121
rect 889 -151 949 -121
rect 979 2230 1009 2379
rect 979 2144 1009 2200
rect 1009 2114 1010 2144
rect 979 2062 1009 2114
rect 979 1944 1009 2032
rect 979 1812 1009 1914
rect 979 1765 1009 1782
rect 1094 1790 1116 1799
rect 1121 1790 1122 1799
rect 1127 1790 1128 1799
rect 1133 1790 1143 1799
rect 1148 1790 1149 1799
rect 1154 1790 1155 1799
rect 1094 1789 1155 1790
rect 1094 1735 1160 1789
rect 979 1562 1009 1735
rect 979 1443 1009 1532
rect 979 1312 1009 1413
rect 979 1214 1009 1282
rect 979 1062 1009 1184
rect 1093 1137 1116 1146
rect 1121 1137 1122 1146
rect 1127 1137 1128 1146
rect 1133 1137 1143 1146
rect 1148 1137 1149 1146
rect 1154 1137 1155 1146
rect 1093 1136 1155 1137
rect 1093 1082 1160 1136
rect 979 812 1009 1032
rect 979 680 1009 782
rect 979 603 1009 650
rect 1009 589 1025 596
rect 1106 645 1125 654
rect 1130 645 1131 654
rect 1136 645 1137 654
rect 1142 645 1152 654
rect 1157 645 1158 654
rect 1163 645 1164 654
rect 1106 644 1164 645
rect 1106 590 1169 644
rect 979 475 1009 573
rect 1009 461 1056 475
rect 979 376 1009 461
rect 1019 460 1056 461
rect 1072 460 1078 475
rect 1619 409 1639 418
rect 1644 409 1645 418
rect 1650 409 1651 418
rect 1656 409 1666 418
rect 1671 409 1672 418
rect 1677 409 1678 418
rect 1619 408 1678 409
rect 1619 354 1683 408
rect 979 321 1009 346
rect 979 218 1009 291
rect 979 214 1059 218
rect 1027 211 1059 214
rect 1068 211 1069 218
rect 979 131 1009 184
rect 1616 155 1636 164
rect 1641 155 1642 164
rect 1647 155 1648 164
rect 1653 155 1663 164
rect 1668 155 1669 164
rect 1674 155 1675 164
rect 1616 154 1675 155
rect 979 31 1009 101
rect 1616 100 1680 154
rect 979 -181 1009 1
rect -1751 -211 -1660 -181
rect -1630 -211 -1540 -181
rect -1510 -211 -1420 -181
rect -1390 -211 -1379 -181
rect -1365 -211 -1300 -181
rect -1270 -211 -1207 -181
rect -1177 -211 -1160 -181
rect -1146 -211 -1060 -181
rect -1030 -211 -940 -181
rect -910 -211 -820 -181
rect -790 -211 -700 -181
rect -670 -211 -580 -181
rect -550 -211 -460 -181
rect -430 -211 -340 -181
rect -310 -211 -220 -181
rect -190 -211 -122 -181
rect -92 -211 -2 -181
rect 28 -211 128 -181
rect 158 -211 248 -181
rect 278 -211 700 -181
rect 730 -211 918 -181
rect 948 -211 1009 -181
rect -1379 -215 -1365 -211
rect -1379 -216 -1317 -215
rect -1160 -216 -1146 -211
rect -1379 -224 -1326 -216
rect -1160 -225 -1124 -216
rect 184 -232 191 -211
rect -945 -285 -881 -266
rect -945 -290 -890 -285
rect -945 -291 -881 -290
rect -945 -296 -890 -291
rect -945 -297 -881 -296
rect -945 -302 -890 -297
rect -945 -312 -881 -302
rect -945 -317 -890 -312
rect -945 -318 -881 -317
rect -945 -323 -890 -318
rect -945 -324 -881 -323
rect -945 -329 -891 -324
rect -446 -285 -382 -266
rect -446 -290 -391 -285
rect -446 -291 -382 -290
rect -446 -296 -391 -291
rect -446 -297 -382 -296
rect -446 -302 -391 -297
rect -446 -312 -382 -302
rect -446 -317 -391 -312
rect -446 -318 -382 -317
rect -446 -323 -391 -318
rect -446 -324 -382 -323
rect -446 -329 -392 -324
rect 185 -332 249 -313
rect 185 -337 240 -332
rect 185 -338 249 -337
rect 185 -343 240 -338
rect 185 -344 249 -343
rect 185 -349 240 -344
rect 185 -359 249 -349
rect 185 -364 240 -359
rect 185 -365 249 -364
rect 185 -370 240 -365
rect 185 -371 249 -370
rect 185 -376 239 -371
rect -1431 -782 -1367 -762
rect -1431 -787 -1376 -782
rect -1431 -788 -1367 -787
rect -1431 -793 -1376 -788
rect -1431 -794 -1367 -793
rect -1431 -799 -1376 -794
rect -1431 -809 -1367 -799
rect -1431 -814 -1376 -809
rect -1431 -815 -1367 -814
rect -1431 -820 -1376 -815
rect -1431 -821 -1367 -820
rect -1431 -826 -1377 -821
rect -1227 -781 -1163 -761
rect -1227 -786 -1172 -781
rect -1227 -787 -1163 -786
rect -1227 -792 -1172 -787
rect -1227 -793 -1163 -792
rect -1227 -798 -1172 -793
rect -1227 -808 -1163 -798
rect -1227 -813 -1172 -808
rect -1227 -814 -1163 -813
rect -1227 -819 -1172 -814
rect -1227 -820 -1163 -819
rect -1227 -825 -1173 -820
<< m234contact >>
rect -1506 3035 -1497 3040
rect -1506 3008 -1497 3013
rect -1291 3035 -1282 3040
rect -1291 3008 -1282 3013
rect -1038 2561 -1029 2566
rect -1038 2534 -1029 2539
rect -791 2561 -782 2566
rect -791 2534 -782 2539
rect -573 2563 -564 2568
rect -573 2536 -564 2541
rect -299 2564 -290 2569
rect -299 2537 -290 2542
rect -1661 2379 -1631 2409
rect -1421 2379 -1391 2409
rect -1181 2379 -1151 2409
rect -941 2379 -911 2409
rect -701 2379 -671 2409
rect -461 2379 -431 2409
rect -221 2379 -191 2409
rect 0 2379 30 2409
rect 207 2379 237 2409
rect 427 2379 457 2409
rect 819 2379 849 2409
rect -1781 2259 -1751 2289
rect -2399 2042 -2394 2051
rect -2372 2042 -2367 2051
rect -1928 1838 -1923 1847
rect -1901 1838 -1896 1847
rect -1781 1779 -1751 1809
rect -1928 1673 -1923 1682
rect -1901 1673 -1896 1682
rect -1929 1438 -1924 1447
rect -1902 1438 -1897 1447
rect -1781 1289 -1751 1319
rect -1929 1181 -1924 1190
rect -1902 1181 -1897 1190
rect -1929 887 -1924 896
rect -1902 887 -1897 896
rect -1781 809 -1751 839
rect -2397 641 -2392 650
rect -2370 641 -2365 650
rect -2397 325 -2392 334
rect -2370 325 -2365 334
rect -1781 339 -1751 369
rect -1781 59 -1751 89
rect -1781 -105 -1751 -75
rect -1721 2319 -1691 2349
rect -1511 2319 -1481 2349
rect -1297 2319 -1267 2349
rect -848 2319 -818 2349
rect -551 2319 -521 2349
rect -311 2319 -281 2349
rect -62 2319 -32 2349
rect 138 2319 168 2349
rect 431 2319 461 2349
rect 729 2319 759 2349
rect -1721 1629 -1691 1659
rect -1721 1139 -1691 1169
rect -1721 659 -1691 689
rect -1721 189 -1691 219
rect -1721 -63 -1691 -33
rect -1601 2259 -1571 2289
rect -1361 2259 -1331 2289
rect -1121 2259 -1091 2289
rect -881 2259 -851 2289
rect -641 2259 -611 2289
rect -401 2259 -371 2289
rect -132 2259 -102 2289
rect 54 2259 84 2289
rect 377 2259 407 2289
rect 642 2259 669 2289
rect -1661 2199 -1631 2229
rect -1661 1719 -1631 1749
rect -1661 1264 -1631 1294
rect -1661 749 -1631 779
rect -1661 279 -1631 309
rect -1661 -1 -1631 29
rect -1451 2199 -1421 2229
rect -1211 2199 -1181 2229
rect -971 2199 -941 2229
rect -731 2199 -701 2229
rect -491 2199 -461 2229
rect -221 2199 -191 2229
rect -6 2199 24 2229
rect 259 2199 289 2229
rect 559 2199 589 2229
rect 789 2199 819 2229
rect -1601 1569 -1571 1599
rect -1601 1079 -1571 1109
rect -1601 599 -1571 629
rect 799 2039 829 2069
rect 799 1880 829 1910
rect 799 1581 829 1611
rect 799 1314 829 1344
rect 799 1085 829 1115
rect 799 601 829 631
rect -1601 129 -1571 159
rect -1450 -31 -1420 -1
rect -1210 -31 -1180 -1
rect -970 -31 -940 -1
rect -730 -31 -700 -1
rect -490 -31 -460 -1
rect -250 -31 -220 -1
rect -32 -31 -2 -1
rect 218 -31 248 -1
rect 790 -31 820 -1
rect 859 2140 889 2170
rect 859 1972 889 2002
rect 859 1722 889 1752
rect 859 1472 889 1502
rect 859 1222 889 1252
rect 859 972 889 1002
rect 859 722 889 752
rect 859 513 889 543
rect 859 231 889 261
rect 859 41 889 71
rect -1599 -91 -1569 -61
rect -1359 -91 -1329 -61
rect -1119 -91 -1089 -61
rect -879 -91 -849 -61
rect -639 -91 -609 -61
rect 59 -91 89 -61
rect 309 -91 339 -61
rect 642 -91 671 -61
rect 919 2118 949 2148
rect 919 1655 949 1685
rect 919 1384 949 1414
rect 919 1152 949 1182
rect 919 594 949 624
rect 919 437 949 467
rect 919 -62 949 -32
rect -1510 -151 -1480 -121
rect -1270 -151 -1240 -121
rect -1030 -151 -1000 -121
rect -790 -151 -760 -121
rect -550 -151 -520 -121
rect -310 -151 -280 -121
rect -92 -151 -62 -121
rect 158 -151 188 -121
rect 730 -151 760 -121
rect 979 2200 1009 2230
rect 979 2032 1009 2062
rect 979 1782 1009 1812
rect 1122 1790 1127 1799
rect 1149 1790 1154 1799
rect 979 1532 1009 1562
rect 979 1282 1009 1312
rect 1122 1137 1127 1146
rect 1149 1137 1154 1146
rect 979 1032 1009 1062
rect 979 782 1009 812
rect 979 573 1009 603
rect 1131 645 1136 654
rect 1158 645 1163 654
rect 1645 409 1650 418
rect 1672 409 1677 418
rect 979 291 1009 321
rect 979 101 1009 131
rect 1642 155 1647 164
rect 1669 155 1674 164
rect -1660 -211 -1630 -181
rect -1420 -211 -1390 -181
rect -1207 -211 -1177 -181
rect -940 -211 -910 -181
rect -700 -211 -670 -181
rect -460 -211 -430 -181
rect -220 -211 -190 -181
rect -2 -211 28 -181
rect 248 -211 278 -181
rect 918 -211 948 -181
rect -890 -296 -881 -291
rect -890 -323 -881 -318
rect -391 -296 -382 -291
rect -391 -323 -382 -318
rect 240 -343 249 -338
rect 240 -370 249 -365
rect -1376 -793 -1367 -788
rect -1376 -820 -1367 -815
rect -1172 -792 -1163 -787
rect -1172 -819 -1163 -814
<< m4contact >>
rect -1721 2055 -1691 2068
rect 919 2067 949 2080
<< metal4 >>
rect -1506 3040 -1442 3046
rect -1497 3035 -1442 3040
rect -1506 3034 -1442 3035
rect -1497 3029 -1442 3034
rect -1506 3028 -1442 3029
rect -1497 3020 -1442 3028
rect -1506 3013 -1442 3020
rect -1497 3008 -1442 3013
rect -1506 3007 -1442 3008
rect -1497 3002 -1442 3007
rect -1506 3001 -1442 3002
rect -1497 2993 -1442 3001
rect -1506 2990 -1442 2993
rect -1291 3040 -1227 3046
rect -1282 3035 -1227 3040
rect -1291 3034 -1227 3035
rect -1282 3029 -1227 3034
rect -1291 3028 -1227 3029
rect -1282 3020 -1227 3028
rect -1291 3013 -1227 3020
rect -1282 3008 -1227 3013
rect -1291 3007 -1227 3008
rect -1282 3002 -1227 3007
rect -1291 3001 -1227 3002
rect -1282 2993 -1227 3001
rect -1291 2990 -1227 2993
rect -1038 2566 -974 2572
rect -1029 2561 -974 2566
rect -1038 2560 -974 2561
rect -1029 2555 -974 2560
rect -1038 2554 -974 2555
rect -1029 2546 -974 2554
rect -1038 2539 -974 2546
rect -1029 2534 -974 2539
rect -1038 2533 -974 2534
rect -1029 2528 -974 2533
rect -1038 2527 -974 2528
rect -1029 2519 -974 2527
rect -1038 2517 -974 2519
rect -791 2566 -727 2572
rect -782 2561 -727 2566
rect -791 2560 -727 2561
rect -782 2555 -727 2560
rect -791 2554 -727 2555
rect -782 2546 -727 2554
rect -791 2539 -727 2546
rect -782 2534 -727 2539
rect -791 2533 -727 2534
rect -782 2528 -727 2533
rect -791 2527 -727 2528
rect -782 2519 -727 2527
rect -791 2517 -727 2519
rect -573 2568 -509 2574
rect -564 2563 -509 2568
rect -573 2562 -509 2563
rect -564 2557 -509 2562
rect -573 2556 -509 2557
rect -564 2548 -509 2556
rect -573 2541 -509 2548
rect -564 2536 -509 2541
rect -573 2535 -509 2536
rect -564 2530 -509 2535
rect -573 2529 -509 2530
rect -564 2521 -509 2529
rect -573 2518 -509 2521
rect -299 2569 -235 2575
rect -290 2564 -235 2569
rect -299 2563 -235 2564
rect -290 2558 -235 2563
rect -299 2557 -235 2558
rect -290 2549 -235 2557
rect -299 2542 -235 2549
rect -290 2537 -235 2542
rect -299 2536 -235 2537
rect -290 2531 -235 2536
rect -299 2530 -235 2531
rect -290 2522 -235 2530
rect -299 2519 -235 2522
rect -1781 2379 -1661 2409
rect -1631 2379 -1421 2409
rect -1391 2379 -1181 2409
rect -1151 2379 -941 2409
rect -911 2379 -701 2409
rect -671 2407 -461 2409
rect -671 2380 -542 2407
rect -513 2380 -461 2407
rect -671 2379 -461 2380
rect -431 2379 -221 2409
rect -191 2379 0 2409
rect 30 2379 207 2409
rect 237 2379 427 2409
rect 457 2379 819 2409
rect 849 2379 1009 2409
rect -1781 2289 -1751 2379
rect -544 2378 -515 2379
rect -269 2349 -240 2351
rect -2405 2051 -2349 2106
rect -2405 2042 -2399 2051
rect -2394 2042 -2393 2051
rect -2388 2042 -2387 2051
rect -2379 2042 -2372 2051
rect -2367 2042 -2366 2051
rect -2361 2042 -2360 2051
rect -2352 2042 -2349 2051
rect -1934 1847 -1879 1902
rect -1934 1838 -1928 1847
rect -1923 1838 -1922 1847
rect -1917 1838 -1916 1847
rect -1908 1838 -1901 1847
rect -1896 1838 -1895 1847
rect -1890 1838 -1889 1847
rect -1881 1838 -1879 1847
rect -1781 1809 -1751 2259
rect -1934 1682 -1879 1737
rect -1934 1673 -1928 1682
rect -1923 1673 -1922 1682
rect -1917 1673 -1916 1682
rect -1908 1673 -1901 1682
rect -1896 1673 -1895 1682
rect -1890 1673 -1889 1682
rect -1881 1673 -1879 1682
rect -1935 1447 -1880 1502
rect -1935 1438 -1929 1447
rect -1924 1438 -1923 1447
rect -1918 1438 -1917 1447
rect -1909 1438 -1902 1447
rect -1897 1438 -1896 1447
rect -1891 1438 -1890 1447
rect -1882 1438 -1880 1447
rect -1781 1319 -1751 1779
rect -1935 1190 -1880 1245
rect -1935 1181 -1929 1190
rect -1924 1181 -1923 1190
rect -1918 1181 -1917 1190
rect -1909 1181 -1902 1190
rect -1897 1181 -1896 1190
rect -1891 1181 -1890 1190
rect -1882 1181 -1880 1190
rect -1935 896 -1880 951
rect -1935 887 -1929 896
rect -1924 887 -1923 896
rect -1918 887 -1917 896
rect -1909 887 -1902 896
rect -1897 887 -1896 896
rect -1891 887 -1890 896
rect -1882 887 -1880 896
rect -1781 839 -1751 1289
rect -2403 650 -2347 705
rect -2403 641 -2397 650
rect -2392 641 -2391 650
rect -2386 641 -2385 650
rect -2377 641 -2370 650
rect -2365 641 -2364 650
rect -2359 641 -2358 650
rect -2350 641 -2347 650
rect -2403 334 -2347 389
rect -2403 325 -2397 334
rect -2392 325 -2391 334
rect -2386 325 -2385 334
rect -2377 325 -2370 334
rect -2365 325 -2364 334
rect -2359 325 -2358 334
rect -2350 325 -2347 334
rect -1781 369 -1751 809
rect -1781 89 -1751 339
rect -1781 -75 -1751 59
rect -1781 -181 -1751 -105
rect -1691 2319 -1511 2349
rect -1481 2319 -1453 2349
rect -1439 2319 -1297 2349
rect -1267 2319 -1246 2349
rect -1216 2319 -1039 2349
rect -1023 2319 -848 2349
rect -818 2319 -792 2349
rect -776 2319 -551 2349
rect -521 2319 -311 2349
rect -281 2348 -62 2349
rect -281 2321 -266 2348
rect -237 2321 -62 2348
rect -281 2319 -62 2321
rect -32 2319 138 2349
rect 168 2319 431 2349
rect 461 2319 729 2349
rect 759 2319 949 2349
rect -1721 2146 -1691 2319
rect -1661 2259 -1601 2289
rect -1571 2259 -1361 2289
rect -1331 2259 -1121 2289
rect -1091 2259 -881 2289
rect -851 2259 -641 2289
rect -611 2259 -557 2289
rect -527 2259 -401 2289
rect -371 2259 -132 2289
rect -102 2259 54 2289
rect 84 2259 377 2289
rect 407 2259 642 2289
rect 669 2259 889 2289
rect -1661 2229 -1631 2259
rect 799 2229 829 2230
rect -1721 2068 -1691 2132
rect -1721 1851 -1691 2055
rect -1721 1686 -1691 1839
rect -1721 1659 -1691 1674
rect -1721 1169 -1691 1629
rect -1721 900 -1691 1139
rect -1721 705 -1691 888
rect -1721 689 -1691 697
rect -1721 389 -1691 659
rect -1721 219 -1691 381
rect -1721 -33 -1691 189
rect -1721 -121 -1691 -63
rect -1661 1749 -1631 2199
rect -1661 1294 -1631 1719
rect -1661 1228 -1631 1264
rect -1661 779 -1631 1198
rect -1661 309 -1631 749
rect -1661 29 -1631 279
rect -1661 -61 -1631 -1
rect -1601 2199 -1451 2229
rect -1421 2199 -1211 2229
rect -1181 2199 -971 2229
rect -941 2199 -731 2229
rect -701 2199 -491 2229
rect -461 2199 -282 2229
rect -252 2199 -221 2229
rect -191 2199 -6 2229
rect 24 2199 259 2229
rect 289 2199 559 2229
rect 589 2199 789 2229
rect 819 2199 829 2229
rect -1601 1599 -1571 2199
rect -1601 1485 -1571 1569
rect -1601 1109 -1571 1455
rect -1601 629 -1571 1079
rect 799 2069 829 2199
rect 799 1910 829 2039
rect 799 1611 829 1880
rect 799 1344 829 1581
rect 799 1115 829 1314
rect 799 631 829 1085
rect -1601 159 -1571 599
rect -1601 -1 -1571 129
rect -1601 -31 -1450 -1
rect -1420 -30 -1314 -1
rect -1306 -2 -1210 -1
rect -1306 -30 -1237 -2
rect -1420 -31 -1237 -30
rect -1229 -31 -1210 -2
rect -1180 -31 -1160 -1
rect -1152 -31 -1085 -1
rect -1077 -31 -1010 -1
rect -1002 -31 -970 -1
rect -940 -31 -928 -1
rect -898 -30 -856 -1
rect -848 -30 -779 -1
rect -898 -31 -779 -30
rect 799 -1 829 601
rect -771 -31 -730 -1
rect -700 -31 -490 -1
rect -460 -31 -250 -1
rect -220 -31 -32 -1
rect -2 -31 218 -1
rect 248 -31 261 -1
rect 274 -31 790 -1
rect 820 -31 829 -1
rect 859 2170 889 2259
rect 859 2002 889 2140
rect 859 1752 889 1972
rect 859 1502 889 1722
rect 859 1252 889 1472
rect 859 1002 889 1222
rect 859 752 889 972
rect 859 543 889 722
rect 859 261 889 513
rect 859 71 889 231
rect -1661 -91 -1599 -61
rect -1569 -91 -1359 -61
rect -1329 -91 -1257 -61
rect -1250 -90 -1180 -61
rect -1173 -90 -1119 -61
rect -1250 -91 -1119 -90
rect -1089 -91 -1029 -61
rect -1022 -91 -879 -61
rect -849 -91 -799 -61
rect -792 -91 -723 -61
rect -716 -91 -639 -61
rect -609 -91 -429 -61
rect -399 -91 59 -61
rect 89 -91 175 -61
rect 859 -61 889 41
rect 186 -91 309 -61
rect 339 -91 642 -61
rect 671 -91 889 -61
rect 919 2148 949 2319
rect 919 2080 949 2118
rect 919 1685 949 2067
rect 919 1414 949 1655
rect 919 1182 949 1384
rect 919 1130 949 1152
rect 919 662 949 1100
rect 919 624 949 632
rect 919 467 949 594
rect 919 420 949 437
rect 919 151 949 407
rect 919 -32 949 138
rect 919 -121 949 -62
rect -1721 -151 -1510 -121
rect -1480 -151 -1433 -121
rect -1420 -151 -1270 -121
rect -1240 -151 -1214 -121
rect -1201 -151 -1030 -121
rect -1000 -151 -790 -121
rect -760 -151 -550 -121
rect -520 -151 -310 -121
rect -280 -151 -92 -121
rect -62 -151 158 -121
rect 188 -150 236 -121
rect 246 -150 730 -121
rect 188 -151 730 -150
rect 760 -151 949 -121
rect 979 2230 1009 2379
rect 979 2062 1009 2200
rect 979 1812 1009 2032
rect 979 1765 1009 1782
rect 1104 1790 1107 1799
rect 1115 1790 1116 1799
rect 1121 1790 1122 1799
rect 1127 1790 1134 1799
rect 1142 1790 1143 1799
rect 1148 1790 1149 1799
rect 1154 1790 1160 1799
rect 1104 1735 1160 1790
rect 979 1562 1009 1735
rect 979 1312 1009 1532
rect 979 1062 1009 1282
rect 1103 1137 1107 1146
rect 1115 1137 1116 1146
rect 1121 1137 1122 1146
rect 1127 1137 1134 1146
rect 1142 1137 1143 1146
rect 1148 1137 1149 1146
rect 1154 1137 1160 1146
rect 1103 1082 1160 1137
rect 979 812 1009 1032
rect 979 603 1009 782
rect 1114 645 1116 654
rect 1124 645 1125 654
rect 1130 645 1131 654
rect 1136 645 1143 654
rect 1151 645 1152 654
rect 1157 645 1158 654
rect 1163 645 1169 654
rect 1114 590 1169 645
rect 979 321 1009 573
rect 1627 409 1630 418
rect 1638 409 1639 418
rect 1644 409 1645 418
rect 1650 409 1657 418
rect 1665 409 1666 418
rect 1671 409 1672 418
rect 1677 409 1683 418
rect 1627 354 1683 409
rect 979 214 1009 291
rect 979 184 1027 214
rect 979 131 1009 184
rect 979 -181 1009 101
rect 1624 155 1627 164
rect 1635 155 1636 164
rect 1641 155 1642 164
rect 1647 155 1654 164
rect 1662 155 1663 164
rect 1668 155 1669 164
rect 1674 155 1680 164
rect 1624 100 1680 155
rect -1781 -211 -1660 -181
rect -1630 -211 -1420 -181
rect -1390 -211 -1207 -181
rect -1177 -211 -940 -181
rect -910 -211 -700 -181
rect -670 -211 -460 -181
rect -430 -211 -220 -181
rect -190 -211 -2 -181
rect 28 -211 248 -181
rect 278 -211 918 -181
rect 948 -211 1009 -181
rect -945 -276 -881 -274
rect -945 -284 -890 -276
rect -945 -285 -881 -284
rect -945 -290 -890 -285
rect -945 -291 -881 -290
rect -945 -296 -890 -291
rect -945 -303 -881 -296
rect -945 -311 -890 -303
rect -945 -312 -881 -311
rect -945 -317 -890 -312
rect -945 -318 -881 -317
rect -945 -323 -890 -318
rect -945 -329 -881 -323
rect -446 -276 -382 -274
rect -446 -284 -391 -276
rect -446 -285 -382 -284
rect -446 -290 -391 -285
rect -446 -291 -382 -290
rect -446 -296 -391 -291
rect -446 -303 -382 -296
rect -446 -311 -391 -303
rect -446 -312 -382 -311
rect -446 -317 -391 -312
rect -446 -318 -382 -317
rect -446 -323 -391 -318
rect -446 -329 -382 -323
rect 185 -323 249 -321
rect 185 -331 240 -323
rect 185 -332 249 -331
rect 185 -337 240 -332
rect 185 -338 249 -337
rect 185 -343 240 -338
rect 185 -350 249 -343
rect 185 -358 240 -350
rect 185 -359 249 -358
rect 185 -364 240 -359
rect 185 -365 249 -364
rect 185 -370 240 -365
rect 185 -376 249 -370
rect -1431 -773 -1367 -770
rect -1431 -781 -1376 -773
rect -1431 -782 -1367 -781
rect -1431 -787 -1376 -782
rect -1431 -788 -1367 -787
rect -1431 -793 -1376 -788
rect -1431 -800 -1367 -793
rect -1431 -808 -1376 -800
rect -1431 -809 -1367 -808
rect -1431 -814 -1376 -809
rect -1431 -815 -1367 -814
rect -1431 -820 -1376 -815
rect -1431 -826 -1367 -820
rect -1227 -772 -1163 -769
rect -1227 -780 -1172 -772
rect -1227 -781 -1163 -780
rect -1227 -786 -1172 -781
rect -1227 -787 -1163 -786
rect -1227 -792 -1172 -787
rect -1227 -799 -1163 -792
rect -1227 -807 -1172 -799
rect -1227 -808 -1163 -807
rect -1227 -813 -1172 -808
rect -1227 -814 -1163 -813
rect -1227 -819 -1172 -814
rect -1227 -825 -1163 -819
<< m345contact >>
rect -1506 3029 -1497 3034
rect -1506 3002 -1497 3007
rect -1291 3029 -1282 3034
rect -1291 3002 -1282 3007
rect -1504 2972 -1444 2978
rect -1289 2972 -1229 2978
rect -1038 2555 -1029 2560
rect -1038 2528 -1029 2533
rect -791 2555 -782 2560
rect -791 2528 -782 2533
rect -573 2557 -564 2562
rect -573 2530 -564 2535
rect -299 2558 -290 2563
rect -299 2531 -290 2536
rect -1038 2497 -974 2505
rect -791 2497 -727 2505
rect -1487 2420 -1466 2438
rect -1267 2433 -1253 2444
rect -1418 2416 -1408 2429
rect -1201 2413 -1192 2434
rect -1039 2421 -1023 2430
rect -1010 2425 -1001 2432
rect -792 2421 -776 2430
rect -762 2427 -753 2433
rect -1801 2134 -1786 2148
rect -2393 2042 -2388 2051
rect -2366 2042 -2361 2051
rect -2337 2044 -2331 2104
rect -1808 2082 -1798 2093
rect -1922 1838 -1917 1847
rect -1895 1838 -1890 1847
rect -1867 1838 -1859 1902
rect -1796 1868 -1791 1873
rect -1793 1839 -1785 1851
rect -1922 1673 -1917 1682
rect -1895 1673 -1890 1682
rect -1867 1673 -1859 1737
rect -1796 1703 -1791 1708
rect -1793 1674 -1785 1686
rect -1923 1438 -1918 1447
rect -1896 1438 -1891 1447
rect -1923 1181 -1918 1190
rect -1896 1181 -1891 1190
rect -1923 887 -1918 896
rect -1896 887 -1891 896
rect -1868 887 -1860 951
rect -1795 917 -1788 923
rect -1794 888 -1786 900
rect -1800 742 -1792 750
rect -2391 641 -2386 650
rect -2364 641 -2359 650
rect -2335 643 -2329 703
rect -1806 684 -1797 690
rect -1797 410 -1787 420
rect -2391 325 -2386 334
rect -2364 325 -2359 334
rect -2335 327 -2329 387
rect -1804 359 -1795 366
rect -1453 2319 -1439 2349
rect -1246 2319 -1216 2349
rect -1039 2319 -1023 2349
rect -792 2319 -776 2349
rect -557 2259 -527 2289
rect -1721 1839 -1691 1851
rect -1721 1674 -1691 1686
rect -1721 888 -1691 900
rect -1721 697 -1691 705
rect -1721 381 -1691 389
rect -1661 1198 -1631 1228
rect -282 2199 -252 2229
rect -1601 1455 -1571 1485
rect 235 596 242 605
rect -285 544 -278 550
rect -694 503 -686 511
rect -639 501 -632 508
rect -582 496 -572 503
rect -494 500 -488 506
rect -479 501 -472 507
rect -428 502 -420 510
rect -376 499 -367 508
rect -330 502 -321 510
rect -67 495 -60 502
rect -495 410 -490 415
rect -218 412 -206 424
rect -230 287 -218 299
rect -499 279 -491 285
rect 207 240 213 252
rect 243 194 250 202
rect 263 198 273 208
rect -1314 182 -1305 190
rect -1238 182 -1229 190
rect -1255 175 -1248 181
rect -1177 174 -1170 180
rect -1161 176 -1152 184
rect -1085 175 -1077 183
rect -1027 175 -1020 181
rect -1010 175 -1002 183
rect -950 176 -943 182
rect -934 173 -926 181
rect -856 177 -848 185
rect -798 174 -791 180
rect -779 176 -771 184
rect -721 172 -713 179
rect -522 174 -514 180
rect -928 -31 -898 -1
rect -429 -91 -399 -61
rect 919 1100 949 1130
rect 919 632 949 662
rect 919 407 949 420
rect 919 138 949 151
rect -1433 -151 -1420 -121
rect -1214 -151 -1201 -121
rect 979 1735 1009 1765
rect 1116 1790 1121 1799
rect 1143 1790 1148 1799
rect 1116 1137 1121 1146
rect 1143 1137 1148 1146
rect 1018 641 1026 653
rect 1017 617 1027 626
rect 1094 590 1102 654
rect 1125 645 1130 654
rect 1152 645 1157 654
rect 1059 376 1069 387
rect 1609 356 1615 416
rect 1639 409 1644 418
rect 1666 409 1671 418
rect 1026 321 1038 333
rect 1051 131 1059 137
rect 1606 102 1612 162
rect 1636 155 1641 164
rect 1663 155 1668 164
rect 1048 73 1057 80
rect -1454 -229 -1446 -220
rect -1408 -224 -1397 -215
rect -1248 -227 -1238 -219
rect -1198 -232 -1191 -226
rect 212 -234 221 -224
rect 236 -233 248 -225
rect -890 -290 -881 -285
rect -890 -317 -881 -312
rect -391 -290 -382 -285
rect 185 -309 249 -301
rect -391 -317 -382 -312
rect 240 -337 249 -332
rect 240 -364 249 -359
rect -1429 -758 -1369 -752
rect -1225 -757 -1165 -751
rect -1376 -787 -1367 -782
rect -1376 -814 -1367 -809
rect -1172 -786 -1163 -781
rect -1172 -813 -1163 -808
<< m5contact >>
rect -542 2380 -513 2407
rect -266 2321 -237 2348
rect -1721 2132 -1690 2146
rect -1314 -30 -1306 -1
rect -1237 -31 -1229 -2
rect -1160 -32 -1152 -1
rect -1085 -32 -1077 -1
rect -1010 -31 -1002 0
rect -856 -30 -848 1
rect -779 -31 -771 0
rect 261 -31 274 -1
rect -1257 -91 -1250 -59
rect -1180 -90 -1173 -58
rect -1029 -91 -1022 -59
rect -799 -93 -792 -61
rect -723 -91 -716 -59
rect 175 -92 186 -60
rect 236 -150 246 -121
<< metal5 >>
rect -1506 3034 -1442 3046
rect -1497 3029 -1442 3034
rect -1506 3028 -1442 3029
rect -1497 3020 -1442 3028
rect -1506 3007 -1442 3020
rect -1497 3002 -1442 3007
rect -1506 3001 -1442 3002
rect -1497 2993 -1442 3001
rect -1506 2990 -1442 2993
rect -1291 3034 -1227 3046
rect -1282 3029 -1227 3034
rect -1291 3028 -1227 3029
rect -1282 3020 -1227 3028
rect -1291 3007 -1227 3020
rect -1282 3002 -1227 3007
rect -1291 3001 -1227 3002
rect -1282 2993 -1227 3001
rect -1291 2990 -1227 2993
rect -1504 2978 -1444 2982
rect -1289 2978 -1229 2982
rect -1038 2560 -974 2572
rect -1029 2555 -974 2560
rect -1038 2554 -974 2555
rect -1029 2546 -974 2554
rect -1038 2533 -974 2546
rect -1029 2528 -974 2533
rect -1038 2527 -974 2528
rect -1029 2519 -974 2527
rect -1038 2517 -974 2519
rect -1038 2505 -974 2509
rect -791 2560 -727 2572
rect -782 2555 -727 2560
rect -791 2554 -727 2555
rect -782 2546 -727 2554
rect -791 2533 -727 2546
rect -782 2528 -727 2533
rect -791 2527 -727 2528
rect -782 2519 -727 2527
rect -791 2517 -727 2519
rect -791 2505 -727 2509
rect -573 2562 -509 2574
rect -564 2557 -509 2562
rect -573 2556 -509 2557
rect -564 2548 -509 2556
rect -573 2535 -509 2548
rect -564 2530 -509 2535
rect -573 2529 -509 2530
rect -564 2521 -509 2529
rect -573 2518 -509 2521
rect -573 2506 -509 2510
rect -299 2563 -235 2575
rect -290 2558 -235 2563
rect -299 2557 -235 2558
rect -290 2549 -235 2557
rect -299 2536 -235 2549
rect -290 2531 -235 2536
rect -299 2530 -235 2531
rect -290 2522 -235 2530
rect -299 2519 -235 2522
rect -1451 2424 -1418 2428
rect -1786 2146 -1689 2148
rect -1786 2134 -1721 2146
rect -1690 2134 -1689 2146
rect -2405 2051 -2349 2106
rect -2405 2042 -2393 2051
rect -2388 2042 -2387 2051
rect -2379 2042 -2366 2051
rect -2361 2042 -2360 2051
rect -2352 2042 -2349 2051
rect -2341 2044 -2337 2104
rect -1486 2099 -1466 2420
rect -1453 2416 -1418 2424
rect -1453 2415 -1408 2416
rect -1453 2349 -1439 2415
rect -1267 2127 -1254 2433
rect -1238 2413 -1201 2426
rect -1013 2432 -999 2441
rect -1238 2412 -1192 2413
rect -1238 2349 -1224 2412
rect -1039 2349 -1023 2421
rect -1013 2425 -1010 2432
rect -1001 2425 -999 2432
rect -764 2433 -750 2438
rect -1013 2157 -999 2425
rect -792 2349 -776 2421
rect -764 2427 -762 2433
rect -753 2427 -750 2433
rect -764 2185 -750 2427
rect -557 2426 -527 2506
rect -299 2498 -235 2511
rect -557 2407 -526 2426
rect -557 2380 -542 2407
rect -557 2375 -526 2380
rect -557 2289 -527 2375
rect -282 2365 -252 2498
rect -282 2348 -251 2365
rect -282 2321 -266 2348
rect -282 2318 -251 2321
rect -282 2229 -252 2318
rect -764 2165 -750 2166
rect 699 2072 700 2084
rect 686 2063 700 2072
rect -1934 1847 -1879 1902
rect -1934 1838 -1922 1847
rect -1917 1838 -1916 1847
rect -1908 1838 -1895 1847
rect -1890 1838 -1889 1847
rect -1881 1838 -1879 1847
rect -1871 1838 -1867 1902
rect -1785 1839 -1721 1851
rect -1934 1682 -1879 1737
rect -1934 1673 -1922 1682
rect -1917 1673 -1916 1682
rect -1908 1673 -1895 1682
rect -1890 1673 -1889 1682
rect -1881 1673 -1879 1682
rect -1871 1673 -1867 1737
rect -1785 1674 -1721 1686
rect -1935 1447 -1880 1502
rect -1935 1438 -1923 1447
rect -1918 1438 -1917 1447
rect -1909 1438 -1896 1447
rect -1891 1438 -1890 1447
rect -1882 1438 -1880 1447
rect -1872 1485 -1859 1502
rect -1872 1455 -1601 1485
rect -1872 1438 -1859 1455
rect -1563 1379 -1556 1868
rect -1569 1369 -1556 1379
rect -1547 1702 -1546 1713
rect -1935 1190 -1880 1245
rect -1935 1181 -1923 1190
rect -1918 1181 -1917 1190
rect -1909 1181 -1896 1190
rect -1891 1181 -1890 1190
rect -1882 1181 -1880 1190
rect -1872 1228 -1846 1245
rect -1872 1198 -1661 1228
rect -1872 1181 -1846 1198
rect -1935 896 -1880 951
rect -1935 887 -1923 896
rect -1918 887 -1917 896
rect -1909 887 -1896 896
rect -1891 887 -1890 896
rect -1882 887 -1880 896
rect -1872 887 -1868 951
rect -1786 888 -1721 900
rect -1792 742 -1783 750
rect -1791 705 -1783 742
rect -2403 650 -2347 705
rect -2403 641 -2391 650
rect -2386 641 -2385 650
rect -2377 641 -2364 650
rect -2359 641 -2358 650
rect -2350 641 -2347 650
rect -2339 643 -2335 703
rect -1791 697 -1721 705
rect -1569 453 -1562 1369
rect -1799 410 -1797 411
rect -1799 389 -1790 410
rect -2403 334 -2347 389
rect -2403 325 -2391 334
rect -2386 325 -2385 334
rect -2377 325 -2364 334
rect -2359 325 -2358 334
rect -2350 325 -2347 334
rect -2339 327 -2335 387
rect -1799 381 -1721 389
rect -1799 380 -1790 381
rect -1547 265 -1539 1702
rect -1488 1454 -1477 2033
rect -1523 191 -1516 915
rect -1487 739 -1480 1454
rect -1487 684 -1479 739
rect -1506 681 -1496 683
rect -1506 557 -1496 671
rect -1486 631 -1479 684
rect -1487 511 -1479 631
rect -696 625 -693 628
rect 686 620 699 2063
rect 712 1983 725 2111
rect 698 604 699 620
rect 711 604 725 1983
rect -656 554 -646 556
rect -656 508 -646 546
rect -479 509 -468 511
rect -427 510 -415 571
rect -117 570 -67 581
rect -133 569 -67 570
rect -286 550 -278 560
rect -286 544 -285 550
rect -582 508 -572 509
rect -1487 500 -1479 502
rect -656 501 -639 508
rect -584 503 -572 508
rect -479 507 -464 509
rect -584 496 -582 503
rect -584 399 -572 496
rect -510 500 -494 506
rect -472 501 -464 507
rect -420 505 -415 510
rect -330 510 -321 512
rect -1406 25 -1405 31
rect -1433 -218 -1420 -151
rect -1406 -215 -1396 25
rect -1313 -1 -1305 182
rect -1306 -30 -1305 -1
rect -1313 -31 -1305 -30
rect -1257 181 -1249 187
rect -1257 175 -1255 181
rect -1257 -59 -1249 175
rect -1237 -2 -1229 182
rect -1180 180 -1172 187
rect -1180 174 -1177 180
rect -1250 -91 -1249 -59
rect -1180 -58 -1172 174
rect -1160 -1 -1152 176
rect -1029 181 -1021 184
rect -1077 175 -1076 180
rect -1084 -1 -1076 175
rect -1077 -5 -1076 -1
rect -1029 175 -1027 181
rect -952 182 -944 187
rect -1002 175 -1001 180
rect -1173 -90 -1172 -58
rect -1180 -91 -1172 -90
rect -1029 -59 -1021 175
rect -1009 0 -1001 175
rect -1002 -5 -1001 0
rect -952 176 -950 182
rect -1022 -91 -1021 -59
rect -952 -91 -944 176
rect -926 173 -924 181
rect -932 0 -924 173
rect -856 1 -848 177
rect -934 -1 -923 0
rect -934 -31 -928 -1
rect -800 180 -792 187
rect -800 174 -798 180
rect -1029 -94 -1021 -91
rect -1214 -202 -1201 -151
rect -1237 -205 -1201 -202
rect -1446 -229 -1420 -218
rect -1397 -220 -1396 -215
rect -1238 -216 -1201 -205
rect -1238 -227 -1227 -216
rect -1214 -218 -1201 -216
rect -928 -262 -898 -31
rect -800 -61 -792 174
rect -779 0 -771 176
rect -723 179 -715 187
rect -723 172 -721 179
rect -800 -91 -799 -61
rect -723 -59 -715 172
rect -510 37 -504 500
rect -479 19 -468 501
rect -367 499 -366 504
rect -374 482 -366 499
rect -330 444 -321 502
rect -286 181 -278 544
rect 711 484 724 604
rect 732 509 745 2140
rect 752 2006 767 2166
rect 753 1485 766 2006
rect 1074 1765 1094 1799
rect 1009 1735 1094 1765
rect 1104 1790 1107 1799
rect 1115 1790 1116 1799
rect 1121 1790 1134 1799
rect 1142 1790 1143 1799
rect 1148 1790 1160 1799
rect 1104 1735 1160 1790
rect 753 1480 767 1485
rect 754 424 767 1480
rect 1073 1130 1093 1146
rect 949 1100 1093 1130
rect 1073 1082 1093 1100
rect 1103 1137 1107 1146
rect 1115 1137 1116 1146
rect 1121 1137 1134 1146
rect 1142 1137 1143 1146
rect 1148 1137 1160 1146
rect 1103 1082 1160 1137
rect 949 641 1018 653
rect 778 583 790 616
rect 1102 590 1106 654
rect 1114 645 1116 654
rect 1124 645 1125 654
rect 1130 645 1143 654
rect 1151 645 1152 654
rect 1157 645 1169 654
rect 1114 590 1169 645
rect 765 414 767 424
rect 777 301 790 583
rect 1026 420 1038 421
rect 949 407 1038 420
rect 1026 333 1038 407
rect 1615 356 1619 416
rect 1627 409 1630 418
rect 1638 409 1639 418
rect 1644 409 1657 418
rect 1665 409 1666 418
rect 1671 409 1683 418
rect 1627 354 1683 409
rect 175 240 207 252
rect 213 240 215 252
rect -716 -91 -715 -59
rect 175 -60 187 240
rect 261 208 272 209
rect 213 200 243 201
rect -429 -262 -399 -91
rect 186 -92 187 -60
rect 212 194 243 200
rect 261 198 263 208
rect 212 193 249 194
rect 212 -224 221 193
rect 261 -1 272 198
rect 1018 151 1028 152
rect 949 138 1028 151
rect 1018 80 1028 138
rect 1612 102 1616 162
rect 1624 155 1627 164
rect 1635 155 1636 164
rect 1641 155 1654 164
rect 1662 155 1663 164
rect 1668 155 1680 164
rect 1624 100 1680 155
rect 1018 73 1048 80
rect 1057 73 1062 80
rect 246 -150 247 -121
rect 236 -216 247 -150
rect 236 -225 248 -216
rect -945 -266 -881 -262
rect -945 -276 -881 -274
rect -945 -284 -890 -276
rect -945 -285 -881 -284
rect -945 -290 -890 -285
rect -945 -303 -881 -290
rect -945 -311 -890 -303
rect -945 -312 -881 -311
rect -945 -317 -890 -312
rect -945 -329 -881 -317
rect -446 -266 -382 -262
rect -446 -276 -382 -274
rect -446 -284 -391 -276
rect -446 -285 -382 -284
rect -446 -290 -391 -285
rect -446 -303 -382 -290
rect -446 -311 -391 -303
rect -446 -312 -382 -311
rect -446 -317 -391 -312
rect -446 -329 -382 -317
rect 185 -313 249 -309
rect 185 -323 249 -321
rect 185 -331 240 -323
rect 185 -332 249 -331
rect 185 -337 240 -332
rect 185 -350 249 -337
rect 185 -358 240 -350
rect 185 -359 249 -358
rect 185 -364 240 -359
rect 185 -376 249 -364
rect -1429 -762 -1369 -758
rect -1225 -761 -1165 -757
rect -1431 -773 -1367 -770
rect -1431 -781 -1376 -773
rect -1431 -782 -1367 -781
rect -1431 -787 -1376 -782
rect -1431 -800 -1367 -787
rect -1431 -808 -1376 -800
rect -1431 -809 -1367 -808
rect -1431 -814 -1376 -809
rect -1431 -826 -1367 -814
rect -1227 -772 -1163 -769
rect -1227 -780 -1172 -772
rect -1227 -781 -1163 -780
rect -1227 -786 -1172 -781
rect -1227 -799 -1163 -786
rect -1227 -807 -1172 -799
rect -1227 -808 -1163 -807
rect -1227 -813 -1172 -808
rect -1227 -825 -1163 -813
<< m456contact >>
rect -1506 3020 -1497 3028
rect -1506 2993 -1497 3001
rect -1506 2982 -1442 2990
rect -1291 3020 -1282 3028
rect -1291 2993 -1282 3001
rect -1291 2982 -1227 2990
rect -1038 2546 -1029 2554
rect -1038 2519 -1029 2527
rect -1038 2509 -974 2517
rect -791 2546 -782 2554
rect -791 2519 -782 2527
rect -791 2509 -727 2517
rect -573 2548 -564 2556
rect -573 2521 -564 2529
rect -573 2510 -509 2518
rect -299 2549 -290 2557
rect -299 2522 -290 2530
rect -299 2511 -235 2519
rect -2387 2042 -2379 2051
rect -2360 2042 -2352 2051
rect -2349 2042 -2341 2106
rect -1916 1838 -1908 1847
rect -1889 1838 -1881 1847
rect -1879 1838 -1871 1902
rect -1916 1673 -1908 1682
rect -1889 1673 -1881 1682
rect -1879 1673 -1871 1737
rect -1917 1438 -1909 1447
rect -1890 1438 -1882 1447
rect -1880 1438 -1872 1502
rect -1917 1181 -1909 1190
rect -1890 1181 -1882 1190
rect -1880 1181 -1872 1245
rect -1917 887 -1909 896
rect -1890 887 -1882 896
rect -1880 887 -1872 951
rect -2385 641 -2377 650
rect -2358 641 -2350 650
rect -2347 641 -2339 705
rect -2385 325 -2377 334
rect -2358 325 -2350 334
rect -2347 325 -2339 389
rect 1094 1735 1104 1799
rect 1107 1790 1115 1799
rect 1134 1790 1142 1799
rect 1093 1082 1103 1146
rect 1107 1137 1115 1146
rect 1134 1137 1142 1146
rect 1106 590 1114 654
rect 1116 645 1124 654
rect 1143 645 1151 654
rect 1619 354 1627 418
rect 1630 409 1638 418
rect 1657 409 1665 418
rect 1616 100 1624 164
rect 1627 155 1635 164
rect 1654 155 1662 164
rect -945 -274 -881 -266
rect -890 -284 -881 -276
rect -890 -311 -881 -303
rect -446 -274 -382 -266
rect -391 -284 -382 -276
rect -391 -311 -382 -303
rect 185 -321 249 -313
rect 240 -331 249 -323
rect 240 -358 249 -350
rect -1431 -770 -1367 -762
rect -1376 -781 -1367 -773
rect -1376 -808 -1367 -800
rect -1227 -769 -1163 -761
rect -1172 -780 -1163 -772
rect -1172 -807 -1163 -799
<< m6contact >>
rect -764 2166 -744 2185
rect 746 2166 770 2185
rect -1014 2138 -994 2157
rect 730 2140 745 2154
rect -1267 2109 -1249 2127
rect 703 2111 728 2130
rect -1798 2082 -1784 2095
rect -1486 2083 -1464 2099
rect 674 2072 699 2093
rect -1492 2033 -1474 2048
rect -1791 1868 -1782 1880
rect -1563 1868 -1553 1879
rect -1791 1703 -1783 1711
rect -1546 1702 -1538 1714
rect -1788 917 -1780 925
rect -1806 675 -1797 684
rect -1569 442 -1559 453
rect -1795 357 -1786 366
rect -1523 915 -1515 926
rect -1547 253 -1535 265
rect -1506 671 -1496 681
rect -1508 541 -1496 557
rect 223 595 235 606
rect 683 604 698 620
rect -427 571 -415 582
rect -657 546 -646 554
rect -1488 502 -1478 511
rect -702 503 -694 511
rect -138 570 -117 582
rect -67 562 -51 581
rect -585 385 -571 399
rect -1523 182 -1514 191
rect -1405 25 -1392 37
rect -1191 -231 -1182 -222
rect -522 180 -514 190
rect -497 415 -489 423
rect -499 271 -491 279
rect -513 25 -504 37
rect -374 469 -366 482
rect -330 433 -321 444
rect -60 495 -52 503
rect 732 492 745 509
rect 709 471 727 484
rect 778 616 791 630
rect 1007 617 1017 626
rect -206 412 -194 424
rect 752 411 765 424
rect 1050 376 1059 387
rect -218 288 -206 300
rect 777 287 791 301
rect -286 165 -275 181
rect -479 10 -470 19
rect 1051 137 1059 146
<< metal6 >>
rect -1506 3028 -1442 3046
rect -1497 3020 -1442 3028
rect -1506 3001 -1442 3020
rect -1497 2993 -1442 3001
rect -1506 2990 -1442 2993
rect -1291 3028 -1227 3046
rect -1282 3020 -1227 3028
rect -1291 3001 -1227 3020
rect -1282 2993 -1227 3001
rect -1291 2990 -1227 2993
rect -1038 2554 -974 2572
rect -1029 2546 -974 2554
rect -1038 2527 -974 2546
rect -1029 2519 -974 2527
rect -1038 2517 -974 2519
rect -791 2554 -727 2572
rect -782 2546 -727 2554
rect -791 2527 -727 2546
rect -782 2519 -727 2527
rect -791 2517 -727 2519
rect -573 2556 -509 2574
rect -564 2548 -509 2556
rect -573 2529 -509 2548
rect -564 2521 -509 2529
rect -573 2518 -509 2521
rect -299 2557 -235 2575
rect -290 2549 -235 2557
rect -299 2530 -235 2549
rect -290 2522 -235 2530
rect -299 2519 -235 2522
rect -328 2184 746 2185
rect -744 2166 746 2184
rect -760 2165 335 2166
rect -994 2153 82 2156
rect -994 2140 730 2153
rect -994 2138 82 2140
rect -997 2137 82 2138
rect -1267 2131 -191 2132
rect -1267 2130 723 2131
rect -1267 2127 703 2130
rect -1249 2112 703 2127
rect -1249 2109 -11 2112
rect -1087 2108 -11 2109
rect -2405 2051 -2349 2106
rect -2405 2042 -2387 2051
rect -2379 2042 -2360 2051
rect -2352 2042 -2349 2051
rect -1490 2083 -1486 2099
rect -1464 2096 -1418 2099
rect -1464 2093 699 2096
rect -1464 2083 674 2093
rect -1797 2045 -1785 2082
rect -1448 2081 674 2083
rect -1521 2045 -1492 2046
rect -1797 2033 -1492 2045
rect -1474 2033 -1472 2046
rect -1797 2032 -1785 2033
rect -1934 1847 -1879 1902
rect -1934 1838 -1916 1847
rect -1908 1838 -1889 1847
rect -1881 1838 -1879 1847
rect -1801 1868 -1791 1874
rect -1782 1879 -1553 1880
rect -1782 1868 -1563 1879
rect -1934 1682 -1879 1737
rect -1934 1673 -1916 1682
rect -1908 1673 -1889 1682
rect -1881 1673 -1879 1682
rect 1104 1790 1107 1799
rect 1115 1790 1134 1799
rect 1142 1790 1160 1799
rect 1104 1735 1160 1790
rect -1783 1713 -1562 1714
rect -1801 1703 -1791 1708
rect -1783 1702 -1546 1713
rect -1538 1702 -1536 1713
rect -1935 1447 -1880 1502
rect -1935 1438 -1917 1447
rect -1909 1438 -1890 1447
rect -1882 1438 -1880 1447
rect -1935 1190 -1880 1245
rect -1935 1181 -1917 1190
rect -1909 1181 -1890 1190
rect -1882 1181 -1880 1190
rect 1103 1137 1107 1146
rect 1115 1137 1134 1146
rect 1142 1137 1160 1146
rect 1103 1082 1160 1137
rect -1935 896 -1880 951
rect -1935 887 -1917 896
rect -1909 887 -1890 896
rect -1882 887 -1880 896
rect -1801 917 -1788 922
rect -1608 922 -1523 923
rect -1780 917 -1523 922
rect -2403 650 -2347 705
rect -2403 641 -2385 650
rect -2377 641 -2358 650
rect -2350 641 -2347 650
rect -1797 675 -1506 681
rect -1806 672 -1506 675
rect -1496 672 -1495 681
rect 258 613 302 617
rect 258 604 683 613
rect 791 617 1007 626
rect 1017 617 1035 626
rect 791 616 1035 617
rect 778 615 1035 616
rect 258 582 270 604
rect 1114 645 1116 654
rect 1124 645 1143 654
rect 1151 645 1169 654
rect 1114 590 1169 645
rect -415 571 -138 581
rect -423 570 -138 571
rect 52 581 270 582
rect -117 570 -116 581
rect -423 568 -116 570
rect -51 563 270 581
rect -51 562 116 563
rect -67 561 -22 562
rect -1496 554 -722 555
rect -1496 546 -657 554
rect -1496 544 -646 546
rect -1478 503 -702 511
rect -694 503 -678 511
rect 514 507 732 508
rect -52 495 732 507
rect 514 491 608 495
rect -374 482 381 483
rect -366 471 709 482
rect -366 469 727 471
rect -28 468 727 469
rect -1570 443 -1569 452
rect -1559 443 -492 452
rect -325 445 545 446
rect -325 444 660 445
rect 1017 444 1059 445
rect -497 423 -492 443
rect -321 435 1060 444
rect -321 433 660 435
rect 1017 434 1060 435
rect -210 432 660 433
rect -497 411 -492 415
rect -222 412 -206 420
rect -194 412 752 420
rect -222 411 752 412
rect -1392 399 -1376 402
rect -2403 334 -2347 389
rect -2403 325 -2385 334
rect -2377 325 -2358 334
rect -2350 325 -2347 334
rect -1392 388 -585 399
rect -1392 387 -596 388
rect -1392 365 -1376 387
rect -571 388 -558 399
rect 1050 387 1060 434
rect 1059 376 1060 387
rect -1489 364 -1374 365
rect -1786 357 -1374 364
rect -1392 356 -1376 357
rect 1627 409 1630 418
rect 1638 409 1657 418
rect 1665 409 1683 418
rect 1627 354 1683 409
rect -232 290 -218 299
rect -500 279 -493 289
rect 772 299 777 300
rect -206 290 777 299
rect 743 289 777 290
rect -500 271 -499 279
rect -500 265 -493 271
rect -1535 255 -493 265
rect -1514 182 -522 190
rect -514 182 -513 190
rect -275 176 794 179
rect -275 165 1059 176
rect 753 163 1059 165
rect 1051 146 1059 163
rect 1624 155 1627 164
rect 1635 155 1654 164
rect 1662 155 1680 164
rect 1624 100 1680 155
rect -1392 35 -697 36
rect -522 35 -513 36
rect -1392 25 -513 35
rect -1186 10 -479 19
rect -1186 7 -470 10
rect -1186 -211 -1177 7
rect -1190 -215 -1177 -211
rect -1191 -218 -1177 -215
rect -1191 -220 -1181 -218
rect -1191 -222 -1182 -220
rect -945 -276 -881 -274
rect -945 -284 -890 -276
rect -945 -303 -881 -284
rect -945 -311 -890 -303
rect -945 -329 -881 -311
rect -446 -276 -382 -274
rect -446 -284 -391 -276
rect -446 -303 -382 -284
rect -446 -311 -391 -303
rect -446 -329 -382 -311
rect 185 -323 249 -321
rect 185 -331 240 -323
rect 185 -350 249 -331
rect 185 -358 240 -350
rect 185 -376 249 -358
rect -1431 -773 -1367 -770
rect -1431 -781 -1376 -773
rect -1431 -800 -1367 -781
rect -1431 -808 -1376 -800
rect -1431 -826 -1367 -808
rect -1227 -772 -1163 -769
rect -1227 -780 -1172 -772
rect -1227 -799 -1163 -780
rect -1227 -807 -1172 -799
rect -1227 -825 -1163 -807
<< glass >>
rect -1497 2991 -1447 3041
rect -1282 2991 -1232 3041
rect -1029 2517 -979 2567
rect -782 2517 -732 2567
rect -564 2519 -514 2569
rect -290 2520 -240 2570
rect -2400 2051 -2350 2101
rect -1929 1847 -1879 1897
rect 1105 1740 1155 1790
rect -1929 1682 -1879 1732
rect -1930 1447 -1880 1497
rect -1930 1190 -1880 1240
rect 1105 1087 1155 1137
rect -1930 896 -1880 946
rect -2398 650 -2348 700
rect 1114 595 1164 645
rect -2398 334 -2348 384
rect 1628 359 1678 409
rect 1625 105 1675 155
rect -940 -324 -890 -274
rect -441 -324 -391 -274
rect 190 -371 240 -321
rect -1426 -821 -1376 -771
rect -1222 -820 -1172 -770
use outputchain  outputchain_0
timestamp 1481052353
transform 0 -1 -1525 1 0 2496
box -50 -119 465 31
use outputchain  outputchain_8
timestamp 1481052353
transform 0 -1 -1310 1 0 2494
box -50 -119 465 31
use outputchain  outputchain_7
timestamp 1481052353
transform -1 0 -1858 0 -1 2026
box -50 -119 465 31
use outputchain  outputchain_6
timestamp 1481052353
transform -1 0 -1850 0 -1 633
box -50 -119 465 31
use outputchain  outputchain_5
timestamp 1481052353
transform -1 0 -1857 0 -1 301
box -50 -119 465 31
use clkdrive  clkdrive_0
timestamp 1480985955
transform 0 -1 247 1 0 239
box -35 -25 326 32
use outputchain  outputchain_1
timestamp 1481052353
transform 1 0 1120 0 1 440
box -50 -119 465 31
use core  core_0
timestamp 1481054563
transform 1 0 -1472 0 1 90
box 0 0 2171 2053
use outputchain  outputchain_2
timestamp 1481052353
transform 1 0 1112 0 1 189
box -50 -119 465 31
use outputchain  outputchain_3
timestamp 1481052353
transform 0 1 -1345 -1 0 -273
box -50 -119 465 31
use outputchain  outputchain_4
timestamp 1481052353
transform 0 1 -1140 -1 0 -276
box -50 -119 465 31
<< labels >>
rlabel metal6 -539 2545 -539 2545 1 Vdd
rlabel metal6 -269 2544 -269 2544 1 Gnd
rlabel metal6 -1912 928 -1912 928 1 input0
rlabel metal6 -1906 1700 -1906 1700 1 input1
rlabel metal6 -1901 1866 -1901 1866 1 input2
rlabel metal6 1142 616 1142 616 1 clear
rlabel metal6 -763 2542 -763 2542 1 calc_hist
rlabel metal6 -1004 2530 -1004 2530 1 read_out
rlabel metal6 221 -346 221 -346 1 clk_top
rlabel metal6 1654 130 1654 130 1 out_valid
rlabel metal6 1645 398 1645 398 1 out_hist0
rlabel metal6 -1395 -801 -1395 -801 1 out_hist4
rlabel metal6 -1202 -785 -1202 -785 1 out_hist3
rlabel metal6 -2377 366 -2377 366 1 out_hist5
rlabel metal6 -2371 683 -2371 683 1 out_hist6
rlabel metal6 -2373 2082 -2373 2082 1 out_hist7
rlabel metal6 -1251 3025 -1251 3025 1 out_hist1
rlabel metal6 -1469 3023 -1469 3023 1 out_hist2
<< end >>
