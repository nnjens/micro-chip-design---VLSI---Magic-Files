magic
tech scmos
timestamp 1481057006
<< metal6 >>
rect 3689 6694 3749 6699
rect 2735 6689 3749 6694
rect 2735 6663 3754 6689
rect 2735 6584 3755 6663
rect 2736 6560 3755 6584
rect 2736 6502 2845 6560
rect 3699 6555 3721 6560
rect 3898 6535 4114 6608
rect 4165 6077 4204 6103
rect 4404 6076 4456 6123
rect 4642 6093 4660 6120
rect 4908 6086 4927 6119
rect 2745 5651 2830 5671
rect 2745 5628 2831 5651
rect 2745 5582 2830 5628
rect 3269 5412 3303 5438
rect 3273 5272 3304 5275
rect 3267 5250 3304 5272
rect 3267 5244 3297 5250
rect 3268 5013 3291 5041
rect 2768 4249 2829 4855
rect 3263 4474 3286 4502
rect 6801 4488 7028 4492
rect 3269 4464 3286 4474
rect 6796 4411 7028 4488
rect 2768 4232 2831 4249
rect 2768 4189 2829 4232
rect 6325 4169 6336 4179
rect 6796 3947 6910 4411
rect 2792 3936 2828 3937
rect 2768 3575 2838 3936
rect 6815 3913 6851 3947
rect 6805 3641 6869 3729
rect 6805 3560 7032 3641
rect 5403 3221 5416 3222
rect 5393 3201 5416 3221
rect 3974 2780 3998 2783
rect 3778 2771 3802 2773
rect 2822 2661 3810 2771
rect 3966 2763 3998 2780
rect 3953 2690 4103 2763
use ninepF  ninepF_8
timestamp 1085807705
transform -1 0 2747 0 -1 6998
box -52 60 3722 857
use ninepF  ninepF_3
timestamp 1085807705
transform 1 0 4112 0 1 6107
box -52 60 3722 857
use ninepF  ninepF_4
timestamp 1085807705
transform -1 0 2751 0 -1 6100
box -52 60 3722 857
use ninepF  ninepF_5
timestamp 1085807705
transform -1 0 2751 0 -1 5265
box -52 60 3722 857
use ninepF  ninepF_2
timestamp 1085807705
transform 1 0 7015 0 1 3995
box -52 60 3722 857
use ninepF  ninepF_6
timestamp 1085807705
transform -1 0 2784 0 -1 4071
box -52 60 3722 857
use ninepF  ninepF_1
timestamp 1085807705
transform 1 0 7015 0 1 3138
box -52 60 3722 857
use chip  chip_0
timestamp 1481056737
transform 1 0 5185 0 1 3556
box -2405 -826 1683 3046
use ninepF  ninepF_7
timestamp 1085807705
transform -1 0 2818 0 -1 3185
box -52 60 3722 857
use ninepF  ninepF_0
timestamp 1085807705
transform 1 0 4160 0 1 2261
box -52 60 3722 857
<< labels >>
rlabel metal6 3284 5422 3284 5422 1 input2
rlabel metal6 3279 5256 3279 5256 1 input1
rlabel metal6 3274 4484 3274 4484 1 input0
rlabel metal6 6830 3954 6830 3954 1 out_hist0
rlabel metal6 6839 3686 6839 3686 1 out_valid
rlabel metal6 6327 4172 6327 4172 1 clear
rlabel metal6 4916 6101 4916 6101 1 Gnd
rlabel metal6 4646 6101 4646 6101 1 Vdd
rlabel metal6 4422 6098 4422 6098 1 calc_hist
rlabel metal6 4180 6086 4180 6086 1 read_out
rlabel metal6 3934 6581 3934 6581 1 out_hist1
rlabel metal6 3716 6579 3716 6579 1 out_hist2
rlabel metal6 2812 5638 2812 5638 1 out_hist7
rlabel metal6 3283 5422 3283 5422 1 input2
rlabel metal6 3279 5257 3279 5257 1 input1
rlabel metal6 3273 4485 3273 4485 1 input0
rlabel metal6 2814 4239 2814 4239 1 out_hist6
rlabel metal6 2808 3922 2808 3922 1 out_hist5
rlabel metal6 3790 2755 3790 2755 1 out_hist4
rlabel metal6 3983 2771 3983 2771 1 out_hist3
rlabel metal6 5406 3209 5406 3209 1 clk_top
<< end >>
