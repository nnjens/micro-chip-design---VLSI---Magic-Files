magic
tech scmos
timestamp 1480978956
<< metal1 >>
rect 17 272 35 280
rect 754 273 755 280
rect 898 274 904 281
rect 1 260 9 267
rect 53 263 61 268
rect 774 263 782 270
rect 830 53 878 62
rect -1 -39 9 12
rect 80 -3 84 4
rect 183 -6 187 1
rect 286 -8 290 1
rect 389 -7 393 1
rect 492 -7 496 1
rect 595 -6 599 1
rect 698 -6 702 1
rect 24 -27 33 -21
rect 774 -39 782 6
rect 951 5 955 6
rect 801 -6 805 1
rect 872 -37 880 3
rect 951 -7 955 3
rect 1054 -3 1058 2
rect 1157 -3 1161 3
rect 1260 -2 1264 3
rect 1363 -2 1367 2
rect 1466 -2 1470 2
rect 1569 -2 1573 3
rect 897 -27 903 -20
rect 1645 -37 1653 5
rect 1672 -2 1676 3
rect 825 -249 873 -240
rect 0 -346 10 -295
rect 80 -304 84 -300
rect 183 -304 187 -299
rect 286 -305 290 -299
rect 389 -307 393 -300
rect 492 -307 496 -300
rect 595 -307 599 -300
rect 698 -307 702 -300
rect 26 -329 35 -323
rect 774 -340 782 -295
rect 801 -307 805 -300
rect 872 -339 880 -299
rect 951 -307 955 -298
rect 1054 -307 1058 -298
rect 1157 -307 1161 -297
rect 1260 -303 1264 -298
rect 1363 -303 1367 -297
rect 1466 -303 1470 -298
rect 1569 -302 1573 -298
rect 897 -329 903 -322
rect 946 -324 959 -323
rect 1049 -324 1062 -323
rect 1152 -324 1165 -323
rect 1255 -324 1268 -323
rect 1645 -338 1653 -296
rect 1672 -303 1676 -299
rect 827 -549 875 -540
rect 0 -644 9 -593
rect 80 -607 84 -601
rect 183 -606 187 -601
rect 286 -606 290 -602
rect 389 -605 393 -601
rect 492 -606 496 -600
rect 595 -609 599 -600
rect 698 -609 702 -601
rect 24 -630 33 -624
rect 618 -629 635 -624
rect 774 -631 782 -595
rect 801 -609 805 -602
rect 872 -630 880 -599
rect 951 -609 955 -600
rect 1054 -609 1058 -601
rect 1157 -609 1161 -601
rect 1260 -609 1264 -601
rect 1363 -609 1367 -601
rect 1466 -605 1470 -600
rect 1569 -606 1573 -600
rect 898 -629 903 -622
rect 945 -624 958 -623
rect 1048 -624 1061 -623
rect 1151 -624 1164 -623
rect 1254 -624 1267 -623
rect 1357 -624 1370 -623
rect 1460 -624 1473 -623
rect 773 -639 782 -631
rect 871 -639 880 -630
rect 1645 -632 1653 -597
rect 1672 -605 1676 -600
rect 1644 -638 1653 -632
rect 1645 -639 1653 -638
rect 774 -640 782 -639
rect 828 -850 876 -841
rect 79 -907 83 -902
rect 182 -907 186 -902
rect 285 -907 289 -902
rect 388 -907 392 -902
rect 491 -907 495 -902
rect 594 -907 598 -902
rect 697 -907 701 -902
rect 800 -907 804 -902
rect 950 -905 954 -900
rect 1053 -905 1057 -901
rect 1156 -906 1160 -901
rect 1259 -905 1263 -901
rect 1362 -905 1366 -901
rect 1465 -904 1469 -901
rect 1568 -904 1572 -901
rect 1671 -904 1675 -901
<< metal2 >>
rect 79 255 83 282
rect 182 256 186 282
rect 285 257 289 282
rect 388 257 392 282
rect 491 256 495 282
rect 594 257 598 282
rect 697 270 701 282
rect 800 270 804 282
rect 1547 275 1610 280
rect 1547 271 1552 275
rect 1605 271 1610 275
rect 871 270 1552 271
rect 800 266 1552 270
rect 1605 266 1675 271
rect 800 265 876 266
rect 697 256 701 265
rect 800 256 804 265
rect 1568 257 1572 266
rect 1671 258 1675 266
rect 774 36 933 45
rect 94 -4 960 1
rect 946 -22 959 -21
rect 1049 -22 1062 -21
rect 197 -26 1063 -22
rect 197 -27 946 -26
rect 959 -27 1049 -26
rect 1062 -27 1063 -26
rect 79 -45 83 -36
rect 182 -46 186 -36
rect 285 -45 289 -36
rect 388 -44 392 -36
rect 491 -45 495 -36
rect 594 -44 598 -36
rect 697 -44 701 -36
rect 800 -44 804 -36
rect 950 -43 954 -35
rect 1053 -44 1057 -35
rect 1156 -43 1160 -35
rect 1259 -43 1263 -35
rect 1362 -43 1366 -35
rect 1465 -44 1469 -35
rect 1568 -44 1572 -35
rect 1671 -44 1675 -35
rect 774 -265 933 -256
rect 300 -305 1166 -300
rect 946 -324 959 -323
rect 1049 -324 1062 -323
rect 1152 -324 1165 -323
rect 1255 -324 1268 -323
rect 403 -328 1269 -324
rect 403 -329 946 -328
rect 959 -329 1049 -328
rect 1062 -329 1152 -328
rect 1165 -329 1255 -328
rect 1268 -329 1269 -328
rect 79 -346 83 -338
rect 182 -347 186 -338
rect 285 -347 289 -338
rect 388 -347 392 -338
rect 491 -347 495 -338
rect 594 -347 598 -338
rect 697 -347 701 -338
rect 800 -346 804 -338
rect 950 -345 954 -337
rect 1053 -346 1057 -337
rect 1156 -346 1160 -337
rect 1259 -345 1263 -337
rect 1362 -347 1366 -337
rect 1465 -346 1469 -337
rect 1568 -346 1572 -337
rect 1671 -345 1675 -337
rect 774 -567 933 -557
rect 506 -607 1372 -602
rect 945 -624 958 -623
rect 1048 -624 1061 -623
rect 1151 -624 1164 -623
rect 1254 -624 1267 -623
rect 1357 -624 1370 -623
rect 1460 -624 1473 -623
rect 609 -628 1475 -624
rect 609 -629 945 -628
rect 958 -629 1048 -628
rect 1061 -629 1151 -628
rect 1164 -629 1254 -628
rect 1267 -629 1357 -628
rect 1370 -629 1460 -628
rect 1473 -629 1475 -628
rect 78 -646 82 -638
rect 181 -647 185 -638
rect 284 -646 288 -638
rect 387 -648 391 -638
rect 490 -646 494 -638
rect 593 -646 597 -638
rect 696 -646 700 -638
rect 799 -647 803 -638
rect 949 -646 953 -637
rect 1052 -646 1056 -637
rect 1155 -645 1159 -637
rect 1258 -647 1262 -637
rect 1361 -645 1365 -637
rect 1464 -645 1468 -637
rect 1567 -646 1571 -637
rect 1670 -646 1674 -637
rect 773 -867 932 -858
<< m3contact >>
rect 697 265 702 270
rect 1567 266 1572 271
rect 78 238 83 243
rect 181 238 186 243
rect 284 238 289 243
rect 387 238 392 243
rect 490 238 495 243
rect 593 238 598 243
rect 696 238 701 243
rect 799 238 804 243
rect 949 239 954 244
rect 1052 239 1057 244
rect 1155 239 1160 244
rect 1258 239 1263 244
rect 1361 239 1366 244
rect 1464 239 1469 244
rect 1567 239 1572 244
rect 1670 239 1675 244
rect 89 -4 94 1
rect 960 -4 965 1
rect 192 -27 197 -22
rect 1063 -27 1068 -22
rect 79 -36 84 -31
rect 182 -36 187 -31
rect 285 -36 290 -31
rect 388 -36 393 -31
rect 491 -36 496 -31
rect 594 -36 599 -31
rect 697 -36 702 -31
rect 800 -36 805 -31
rect 950 -35 955 -30
rect 1053 -35 1058 -30
rect 1156 -35 1161 -30
rect 1259 -35 1264 -30
rect 1362 -35 1367 -30
rect 1465 -35 1470 -30
rect 1568 -35 1573 -30
rect 1671 -35 1676 -30
rect 78 -63 83 -58
rect 181 -63 186 -58
rect 284 -63 289 -58
rect 387 -63 392 -58
rect 490 -63 495 -58
rect 593 -63 598 -58
rect 696 -63 701 -58
rect 799 -63 804 -58
rect 949 -62 954 -57
rect 1052 -62 1057 -57
rect 1155 -62 1160 -57
rect 1258 -62 1263 -57
rect 1361 -62 1366 -57
rect 1464 -62 1469 -57
rect 1567 -62 1572 -57
rect 1670 -62 1675 -57
rect 295 -305 300 -300
rect 1166 -305 1171 -300
rect 398 -329 403 -324
rect 1269 -329 1274 -324
rect 79 -338 84 -333
rect 182 -338 187 -333
rect 285 -338 290 -333
rect 388 -338 393 -333
rect 491 -338 496 -333
rect 594 -338 599 -333
rect 697 -338 702 -333
rect 800 -338 805 -333
rect 950 -337 955 -332
rect 1053 -337 1058 -332
rect 1156 -337 1161 -332
rect 1259 -337 1264 -332
rect 1362 -337 1367 -332
rect 1465 -337 1470 -332
rect 1568 -337 1573 -332
rect 1671 -337 1676 -332
rect 78 -365 83 -360
rect 181 -365 186 -360
rect 284 -365 289 -360
rect 387 -365 392 -360
rect 490 -365 495 -360
rect 593 -365 598 -360
rect 696 -365 701 -360
rect 799 -365 804 -360
rect 949 -364 954 -359
rect 1052 -364 1057 -359
rect 1155 -364 1160 -359
rect 1258 -364 1263 -359
rect 1361 -364 1366 -359
rect 1464 -364 1469 -359
rect 1567 -364 1572 -359
rect 1670 -364 1675 -359
rect 501 -607 506 -602
rect 1372 -607 1377 -602
rect 604 -629 609 -624
rect 1475 -629 1480 -624
rect 78 -638 83 -633
rect 181 -638 186 -633
rect 284 -638 289 -633
rect 387 -638 392 -633
rect 490 -638 495 -633
rect 593 -638 598 -633
rect 696 -638 701 -633
rect 799 -638 804 -633
rect 949 -637 954 -632
rect 1052 -637 1057 -632
rect 1155 -637 1160 -632
rect 1258 -637 1263 -632
rect 1361 -637 1366 -632
rect 1464 -637 1469 -632
rect 1567 -637 1572 -632
rect 1670 -637 1675 -632
<< m123contact >>
rect 909 -53 914 -48
<< metal3 >>
rect 871 270 1567 271
rect 702 266 1567 270
rect 702 265 876 266
rect -5 256 27 261
rect 886 257 897 262
rect -5 247 43 252
rect 887 248 913 253
rect 83 238 94 243
rect 186 238 197 243
rect 289 238 300 243
rect 392 238 403 243
rect 495 238 506 243
rect 598 238 609 243
rect 701 238 712 243
rect 804 238 815 243
rect 954 239 965 244
rect 1057 239 1068 244
rect 1160 239 1171 244
rect 1263 239 1274 244
rect 1366 239 1377 244
rect 1469 239 1480 244
rect 1572 239 1583 244
rect 1675 239 1686 244
rect 89 1 94 238
rect 89 -31 94 -4
rect 192 -22 197 238
rect 192 -31 197 -27
rect 295 -31 300 238
rect 398 -31 403 238
rect 501 -31 506 238
rect 604 -31 609 238
rect 707 -31 712 238
rect 810 -31 815 238
rect 960 1 965 239
rect 960 -30 965 -4
rect 1063 -22 1068 239
rect 1063 -30 1068 -27
rect 1166 -30 1171 239
rect 1269 -30 1274 239
rect 1372 -30 1377 239
rect 1475 -30 1480 239
rect 1578 -30 1583 239
rect 1681 -30 1686 239
rect 84 -36 94 -31
rect 187 -36 197 -31
rect 290 -36 300 -31
rect 393 -36 403 -31
rect 496 -36 506 -31
rect 599 -36 609 -31
rect 702 -36 712 -31
rect 805 -36 815 -31
rect 955 -35 965 -30
rect 1058 -35 1068 -30
rect 1161 -35 1171 -30
rect 1264 -35 1274 -30
rect 1367 -35 1377 -30
rect 1470 -35 1480 -30
rect 1573 -35 1583 -30
rect 1676 -35 1686 -30
rect 10 -45 27 -40
rect 885 -44 896 -39
rect 10 -54 43 -49
rect 863 -53 909 -48
rect 83 -63 94 -58
rect 186 -63 197 -58
rect 289 -63 300 -58
rect 392 -63 403 -58
rect 495 -63 506 -58
rect 598 -63 609 -58
rect 701 -63 712 -58
rect 804 -63 815 -58
rect 954 -62 965 -57
rect 1057 -62 1068 -57
rect 1160 -62 1171 -57
rect 1263 -62 1274 -57
rect 1366 -61 1377 -57
rect 89 -333 94 -63
rect 192 -333 197 -63
rect 295 -300 300 -63
rect 295 -333 300 -305
rect 398 -324 403 -63
rect 398 -333 403 -329
rect 501 -333 506 -63
rect 604 -333 609 -63
rect 707 -333 712 -63
rect 810 -333 815 -63
rect 960 -332 965 -62
rect 1063 -332 1068 -62
rect 1166 -300 1171 -62
rect 1166 -332 1171 -305
rect 1269 -324 1274 -62
rect 1269 -332 1274 -329
rect 1372 -332 1377 -61
rect 1469 -62 1480 -57
rect 1572 -62 1583 -57
rect 1675 -62 1686 -57
rect 1475 -332 1480 -62
rect 1578 -332 1583 -62
rect 1681 -332 1686 -62
rect 84 -338 94 -333
rect 187 -338 197 -333
rect 290 -338 300 -333
rect 393 -338 403 -333
rect 496 -338 506 -333
rect 599 -338 609 -333
rect 702 -338 712 -333
rect 805 -338 815 -333
rect 955 -337 965 -332
rect 1058 -337 1068 -332
rect 1161 -337 1171 -332
rect 1264 -337 1274 -332
rect 1367 -337 1377 -332
rect 1470 -337 1480 -332
rect 1573 -337 1583 -332
rect 1676 -337 1686 -332
rect 7 -347 27 -342
rect 887 -346 894 -341
rect 7 -356 40 -351
rect 888 -355 913 -350
rect 83 -365 94 -360
rect 186 -365 197 -360
rect 289 -365 300 -360
rect 392 -365 403 -360
rect 495 -365 506 -360
rect 598 -365 609 -360
rect 701 -365 712 -360
rect 804 -365 815 -360
rect 954 -364 965 -359
rect 1057 -364 1068 -359
rect 1160 -364 1171 -359
rect 1263 -364 1274 -359
rect 1366 -364 1377 -359
rect 1469 -364 1480 -359
rect 1572 -364 1583 -359
rect 1675 -364 1686 -359
rect 89 -633 94 -365
rect 192 -633 197 -365
rect 295 -633 300 -365
rect 398 -633 403 -365
rect 501 -602 506 -365
rect 501 -633 506 -607
rect 604 -624 609 -365
rect 604 -633 609 -629
rect 707 -633 712 -365
rect 810 -633 815 -365
rect 960 -632 965 -364
rect 1063 -632 1068 -364
rect 1166 -632 1171 -364
rect 1269 -632 1274 -364
rect 1372 -602 1377 -364
rect 1372 -632 1377 -607
rect 1475 -624 1480 -364
rect 1475 -632 1480 -629
rect 1578 -632 1583 -364
rect 1681 -632 1686 -364
rect 83 -638 94 -633
rect 186 -638 197 -633
rect 289 -638 300 -633
rect 392 -638 403 -633
rect 495 -638 506 -633
rect 598 -638 609 -633
rect 701 -638 712 -633
rect 804 -638 815 -633
rect 954 -637 965 -632
rect 1057 -637 1068 -632
rect 1160 -637 1171 -632
rect 1263 -637 1274 -632
rect 1366 -637 1377 -632
rect 1469 -637 1480 -632
rect 1572 -637 1583 -632
rect 1675 -637 1686 -632
rect -4 -647 24 -642
rect 885 -646 896 -641
rect -5 -656 41 -651
rect 885 -655 912 -650
use word  word_0
timestamp 1480562330
transform 1 0 56 0 1 721
box -56 -721 777 -441
use word  word_4
timestamp 1480562330
transform 1 0 927 0 1 722
box -56 -721 777 -441
use word  word_1
timestamp 1480562330
transform 1 0 56 0 1 420
box -56 -721 777 -441
use word  word_5
timestamp 1480562330
transform 1 0 927 0 1 421
box -56 -721 777 -441
use word  word_2
timestamp 1480562330
transform 1 0 56 0 1 118
box -56 -721 777 -441
use word  word_6
timestamp 1480562330
transform 1 0 927 0 1 119
box -56 -721 777 -441
use word  word_3
timestamp 1480562330
transform 1 0 55 0 1 -182
box -56 -721 777 -441
use word  word_7
timestamp 1480562330
transform 1 0 926 0 1 -181
box -56 -721 777 -441
<< labels >>
rlabel metal2 802 281 802 281 1 new0
rlabel metal1 4 264 4 264 3 Vdd
rlabel metal1 57 266 57 266 1 Gnd
rlabel metal1 22 277 22 277 1 clk0
rlabel metal1 29 -326 29 -326 1 clk2
rlabel metal1 28 -628 28 -628 1 clk3
rlabel metal1 900 278 900 278 1 clk4
rlabel metal1 899 -21 899 -21 1 clk5
rlabel metal1 900 -323 900 -323 1 clk6
rlabel metal1 900 -623 900 -623 1 clk7
rlabel metal3 -3 258 -3 258 3 en0
rlabel metal3 -3 249 -3 249 3 Nen0
rlabel metal1 26 -24 26 -24 1 clk1
rlabel metal3 -3 -645 -3 -645 1 en3
rlabel metal3 -3 -653 -3 -653 1 Nen3
rlabel metal3 888 259 888 259 1 en4
rlabel metal3 890 251 890 251 1 Nen4
rlabel metal3 889 -41 889 -41 1 en5
rlabel metal3 890 -343 890 -343 1 en6
rlabel metal3 891 -353 891 -353 1 Nen6
rlabel metal3 887 -643 887 -643 1 en7
rlabel metal3 888 -652 888 -652 1 Nen7
rlabel metal1 82 -1 82 -1 1 Q0_7
rlabel metal1 185 -5 185 -5 1 Q0_6
rlabel metal1 288 -6 288 -6 1 Q0_5
rlabel metal1 391 -6 391 -6 1 Q0_4
rlabel metal1 494 -5 494 -5 1 Q0_3
rlabel metal1 597 -5 597 -5 1 Q0_2
rlabel metal1 700 -5 700 -5 1 Q0_1
rlabel metal1 803 -5 803 -5 1 Q0_0
rlabel metal1 82 -302 82 -302 1 Q1_7
rlabel metal1 185 -302 185 -302 1 Q1_6
rlabel metal1 288 -303 288 -303 1 Q1_5
rlabel metal1 391 -306 391 -306 1 Q1_4
rlabel metal1 494 -306 494 -306 1 Q1_3
rlabel metal1 597 -306 597 -306 1 Q1_2
rlabel metal1 700 -306 700 -306 1 Q1_1
rlabel metal1 803 -306 803 -306 1 Q1_0
rlabel metal1 82 -605 82 -605 1 Q2_7
rlabel metal1 184 -604 184 -604 1 Q2_6
rlabel metal1 288 -604 288 -604 1 Q2_5
rlabel metal1 391 -603 391 -603 1 Q2_4
rlabel metal1 494 -603 494 -603 1 Q2_3
rlabel metal1 597 -608 597 -608 1 Q2_2
rlabel metal1 700 -608 700 -608 1 Q2_1
rlabel metal1 803 -608 803 -608 1 Q2_0
rlabel metal1 81 -905 81 -905 1 Q3_7
rlabel metal1 184 -905 184 -905 1 Q3_6
rlabel metal1 287 -905 287 -905 1 Q3_5
rlabel metal1 390 -905 390 -905 1 Q3_4
rlabel metal1 493 -905 493 -905 1 Q3_3
rlabel metal1 596 -905 596 -905 1 Q3_2
rlabel metal1 699 -905 699 -905 1 Q3_1
rlabel metal1 802 -905 802 -905 1 Q3_0
rlabel metal1 953 -5 953 -5 1 Q4_7
rlabel metal1 1056 0 1056 0 1 Q4_6
rlabel metal1 1159 -1 1159 -1 1 Q4_5
rlabel metal1 1262 0 1262 0 1 Q4_4
rlabel metal1 1365 -1 1365 -1 1 Q4_3
rlabel metal1 1468 0 1468 0 1 Q4_2
rlabel metal1 1571 0 1571 0 1 Q4_1
rlabel metal1 1674 0 1674 0 1 Q4_0
rlabel metal1 953 -306 953 -306 1 Q5_7
rlabel metal1 1055 -306 1055 -306 1 Q5_6
rlabel metal1 1159 -306 1159 -306 1 Q5_5
rlabel metal1 1262 -301 1262 -301 1 Q5_4
rlabel metal1 1365 -302 1365 -302 1 Q5_3
rlabel metal1 1468 -301 1468 -301 1 Q5_2
rlabel metal1 1572 -301 1572 -301 1 Q5_1
rlabel metal1 1674 -301 1674 -301 1 Q5_0
rlabel metal1 953 -608 953 -608 1 Q6_7
rlabel metal1 1056 -608 1056 -608 1 Q6_6
rlabel metal1 1159 -608 1159 -608 1 Q6_5
rlabel metal1 1262 -608 1262 -608 1 Q6_4
rlabel metal1 1365 -608 1365 -608 1 Q6_3
rlabel metal1 1468 -604 1468 -604 1 Q6_2
rlabel metal1 1571 -604 1571 -604 1 Q6_1
rlabel metal1 1674 -603 1674 -603 1 Q6_0
rlabel metal1 952 -903 952 -903 1 Q7_7
rlabel metal1 1055 -903 1055 -903 1 Q7_6
rlabel metal1 1158 -904 1158 -904 1 Q7_5
rlabel metal1 1261 -903 1261 -903 1 Q7_4
rlabel metal1 1364 -903 1364 -903 1 Q7_3
rlabel metal1 1467 -903 1467 -903 1 Q7_2
rlabel metal1 1570 -903 1570 -903 1 Q7_1
rlabel metal1 1673 -903 1673 -903 1 Q7_0
rlabel metal3 865 -51 865 -51 1 Nen5
rlabel metal2 698 281 698 281 5 new1
rlabel metal2 595 281 595 281 5 new2
rlabel metal2 492 281 492 281 5 new3
rlabel metal2 389 281 389 281 5 new4
rlabel metal2 286 281 286 281 5 new5
rlabel metal2 183 281 183 281 5 new6
rlabel metal2 81 281 81 281 5 new7
rlabel metal3 13 -346 13 -346 1 en2
rlabel metal3 13 -353 13 -353 1 Nen2
rlabel metal3 14 -43 14 -43 1 en1
rlabel metal3 14 -51 14 -51 1 Nen1
<< end >>
