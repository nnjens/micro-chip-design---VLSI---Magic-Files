magic
tech scmos
timestamp 1480976721
<< nwell >>
rect 24 -21 347 20
rect 24 -97 347 -56
rect 24 -173 347 -132
rect 24 -249 347 -208
rect 24 -325 347 -284
rect 24 -401 347 -360
rect 24 -477 347 -436
rect 24 -553 347 -512
<< pwell >>
rect 24 -56 347 -21
rect 24 -126 347 -97
rect 24 -208 347 -173
rect 24 -278 347 -249
rect 24 -360 347 -325
rect 24 -430 347 -401
rect 24 -512 347 -477
rect 24 -582 347 -553
<< ntransistor >>
rect 48 -34 50 -30
rect 60 -34 62 -30
rect 82 -34 84 -30
rect 94 -34 96 -30
rect 116 -34 118 -30
rect 128 -34 130 -30
rect 150 -34 152 -30
rect 162 -34 164 -30
rect 184 -34 186 -30
rect 196 -34 198 -30
rect 218 -34 220 -30
rect 230 -34 232 -30
rect 252 -34 254 -30
rect 264 -34 266 -30
rect 286 -34 288 -30
rect 298 -34 300 -30
rect 320 -34 322 -30
rect 332 -34 334 -30
rect 48 -110 50 -106
rect 60 -110 62 -106
rect 82 -110 84 -106
rect 94 -110 96 -106
rect 116 -110 118 -106
rect 128 -110 130 -106
rect 150 -110 152 -106
rect 162 -110 164 -106
rect 184 -110 186 -106
rect 196 -110 198 -106
rect 218 -110 220 -106
rect 230 -110 232 -106
rect 252 -110 254 -106
rect 264 -110 266 -106
rect 286 -110 288 -106
rect 298 -110 300 -106
rect 320 -110 322 -106
rect 332 -110 334 -106
rect 48 -186 50 -182
rect 60 -186 62 -182
rect 82 -186 84 -182
rect 94 -186 96 -182
rect 116 -186 118 -182
rect 128 -186 130 -182
rect 150 -186 152 -182
rect 162 -186 164 -182
rect 184 -186 186 -182
rect 196 -186 198 -182
rect 218 -186 220 -182
rect 230 -186 232 -182
rect 252 -186 254 -182
rect 264 -186 266 -182
rect 286 -186 288 -182
rect 298 -186 300 -182
rect 320 -186 322 -182
rect 332 -186 334 -182
rect 48 -262 50 -258
rect 60 -262 62 -258
rect 82 -262 84 -258
rect 94 -262 96 -258
rect 116 -262 118 -258
rect 128 -262 130 -258
rect 150 -262 152 -258
rect 162 -262 164 -258
rect 184 -262 186 -258
rect 196 -262 198 -258
rect 218 -262 220 -258
rect 230 -262 232 -258
rect 252 -262 254 -258
rect 264 -262 266 -258
rect 286 -262 288 -258
rect 298 -262 300 -258
rect 320 -262 322 -258
rect 332 -262 334 -258
rect 48 -338 50 -334
rect 60 -338 62 -334
rect 82 -338 84 -334
rect 94 -338 96 -334
rect 116 -338 118 -334
rect 128 -338 130 -334
rect 150 -338 152 -334
rect 162 -338 164 -334
rect 184 -338 186 -334
rect 196 -338 198 -334
rect 218 -338 220 -334
rect 230 -338 232 -334
rect 252 -338 254 -334
rect 264 -338 266 -334
rect 286 -338 288 -334
rect 298 -338 300 -334
rect 320 -338 322 -334
rect 332 -338 334 -334
rect 48 -414 50 -410
rect 60 -414 62 -410
rect 82 -414 84 -410
rect 94 -414 96 -410
rect 116 -414 118 -410
rect 128 -414 130 -410
rect 150 -414 152 -410
rect 162 -414 164 -410
rect 184 -414 186 -410
rect 196 -414 198 -410
rect 218 -414 220 -410
rect 230 -414 232 -410
rect 252 -414 254 -410
rect 264 -414 266 -410
rect 286 -414 288 -410
rect 298 -414 300 -410
rect 320 -414 322 -410
rect 332 -414 334 -410
rect 48 -490 50 -486
rect 60 -490 62 -486
rect 82 -490 84 -486
rect 94 -490 96 -486
rect 116 -490 118 -486
rect 128 -490 130 -486
rect 150 -490 152 -486
rect 162 -490 164 -486
rect 184 -490 186 -486
rect 196 -490 198 -486
rect 218 -490 220 -486
rect 230 -490 232 -486
rect 252 -490 254 -486
rect 264 -490 266 -486
rect 286 -490 288 -486
rect 298 -490 300 -486
rect 320 -490 322 -486
rect 332 -490 334 -486
rect 48 -566 50 -562
rect 60 -566 62 -562
rect 82 -566 84 -562
rect 94 -566 96 -562
rect 116 -566 118 -562
rect 128 -566 130 -562
rect 150 -566 152 -562
rect 162 -566 164 -562
rect 184 -566 186 -562
rect 196 -566 198 -562
rect 218 -566 220 -562
rect 230 -566 232 -562
rect 252 -566 254 -562
rect 264 -566 266 -562
rect 286 -566 288 -562
rect 298 -566 300 -562
rect 320 -566 322 -562
rect 332 -566 334 -562
<< ptransistor >>
rect 48 0 50 6
rect 60 0 62 6
rect 82 0 84 6
rect 94 0 96 6
rect 116 0 118 6
rect 128 0 130 6
rect 150 0 152 6
rect 162 0 164 6
rect 184 0 186 6
rect 196 0 198 6
rect 218 0 220 6
rect 230 0 232 6
rect 252 0 254 6
rect 264 0 266 6
rect 286 0 288 6
rect 298 0 300 6
rect 320 0 322 6
rect 332 0 334 6
rect 48 -76 50 -70
rect 60 -76 62 -70
rect 82 -76 84 -70
rect 94 -76 96 -70
rect 116 -76 118 -70
rect 128 -76 130 -70
rect 150 -76 152 -70
rect 162 -76 164 -70
rect 184 -76 186 -70
rect 196 -76 198 -70
rect 218 -76 220 -70
rect 230 -76 232 -70
rect 252 -76 254 -70
rect 264 -76 266 -70
rect 286 -76 288 -70
rect 298 -76 300 -70
rect 320 -76 322 -70
rect 332 -76 334 -70
rect 48 -152 50 -146
rect 60 -152 62 -146
rect 82 -152 84 -146
rect 94 -152 96 -146
rect 116 -152 118 -146
rect 128 -152 130 -146
rect 150 -152 152 -146
rect 162 -152 164 -146
rect 184 -152 186 -146
rect 196 -152 198 -146
rect 218 -152 220 -146
rect 230 -152 232 -146
rect 252 -152 254 -146
rect 264 -152 266 -146
rect 286 -152 288 -146
rect 298 -152 300 -146
rect 320 -152 322 -146
rect 332 -152 334 -146
rect 48 -228 50 -222
rect 60 -228 62 -222
rect 82 -228 84 -222
rect 94 -228 96 -222
rect 116 -228 118 -222
rect 128 -228 130 -222
rect 150 -228 152 -222
rect 162 -228 164 -222
rect 184 -228 186 -222
rect 196 -228 198 -222
rect 218 -228 220 -222
rect 230 -228 232 -222
rect 252 -228 254 -222
rect 264 -228 266 -222
rect 286 -228 288 -222
rect 298 -228 300 -222
rect 320 -228 322 -222
rect 332 -228 334 -222
rect 48 -304 50 -298
rect 60 -304 62 -298
rect 82 -304 84 -298
rect 94 -304 96 -298
rect 116 -304 118 -298
rect 128 -304 130 -298
rect 150 -304 152 -298
rect 162 -304 164 -298
rect 184 -304 186 -298
rect 196 -304 198 -298
rect 218 -304 220 -298
rect 230 -304 232 -298
rect 252 -304 254 -298
rect 264 -304 266 -298
rect 286 -304 288 -298
rect 298 -304 300 -298
rect 320 -304 322 -298
rect 332 -304 334 -298
rect 48 -380 50 -374
rect 60 -380 62 -374
rect 82 -380 84 -374
rect 94 -380 96 -374
rect 116 -380 118 -374
rect 128 -380 130 -374
rect 150 -380 152 -374
rect 162 -380 164 -374
rect 184 -380 186 -374
rect 196 -380 198 -374
rect 218 -380 220 -374
rect 230 -380 232 -374
rect 252 -380 254 -374
rect 264 -380 266 -374
rect 286 -380 288 -374
rect 298 -380 300 -374
rect 320 -380 322 -374
rect 332 -380 334 -374
rect 48 -456 50 -450
rect 60 -456 62 -450
rect 82 -456 84 -450
rect 94 -456 96 -450
rect 116 -456 118 -450
rect 128 -456 130 -450
rect 150 -456 152 -450
rect 162 -456 164 -450
rect 184 -456 186 -450
rect 196 -456 198 -450
rect 218 -456 220 -450
rect 230 -456 232 -450
rect 252 -456 254 -450
rect 264 -456 266 -450
rect 286 -456 288 -450
rect 298 -456 300 -450
rect 320 -456 322 -450
rect 332 -456 334 -450
rect 48 -532 50 -526
rect 60 -532 62 -526
rect 82 -532 84 -526
rect 94 -532 96 -526
rect 116 -532 118 -526
rect 128 -532 130 -526
rect 150 -532 152 -526
rect 162 -532 164 -526
rect 184 -532 186 -526
rect 196 -532 198 -526
rect 218 -532 220 -526
rect 230 -532 232 -526
rect 252 -532 254 -526
rect 264 -532 266 -526
rect 286 -532 288 -526
rect 298 -532 300 -526
rect 320 -532 322 -526
rect 332 -532 334 -526
<< ndiffusion >>
rect 45 -34 48 -30
rect 50 -34 60 -30
rect 62 -34 65 -30
rect 79 -34 82 -30
rect 84 -34 94 -30
rect 96 -34 99 -30
rect 113 -34 116 -30
rect 118 -34 128 -30
rect 130 -34 133 -30
rect 147 -34 150 -30
rect 152 -34 162 -30
rect 164 -34 167 -30
rect 181 -34 184 -30
rect 186 -34 196 -30
rect 198 -34 201 -30
rect 215 -34 218 -30
rect 220 -34 230 -30
rect 232 -34 235 -30
rect 249 -34 252 -30
rect 254 -34 264 -30
rect 266 -34 269 -30
rect 283 -34 286 -30
rect 288 -34 298 -30
rect 300 -34 303 -30
rect 317 -34 320 -30
rect 322 -34 332 -30
rect 334 -34 337 -30
rect 45 -110 48 -106
rect 50 -110 60 -106
rect 62 -110 65 -106
rect 79 -110 82 -106
rect 84 -110 94 -106
rect 96 -110 99 -106
rect 113 -110 116 -106
rect 118 -110 128 -106
rect 130 -110 133 -106
rect 147 -110 150 -106
rect 152 -110 162 -106
rect 164 -110 167 -106
rect 181 -110 184 -106
rect 186 -110 196 -106
rect 198 -110 201 -106
rect 215 -110 218 -106
rect 220 -110 230 -106
rect 232 -110 235 -106
rect 249 -110 252 -106
rect 254 -110 264 -106
rect 266 -110 269 -106
rect 283 -110 286 -106
rect 288 -110 298 -106
rect 300 -110 303 -106
rect 317 -110 320 -106
rect 322 -110 332 -106
rect 334 -110 337 -106
rect 45 -186 48 -182
rect 50 -186 60 -182
rect 62 -186 65 -182
rect 79 -186 82 -182
rect 84 -186 94 -182
rect 96 -186 99 -182
rect 113 -186 116 -182
rect 118 -186 128 -182
rect 130 -186 133 -182
rect 147 -186 150 -182
rect 152 -186 162 -182
rect 164 -186 167 -182
rect 181 -186 184 -182
rect 186 -186 196 -182
rect 198 -186 201 -182
rect 215 -186 218 -182
rect 220 -186 230 -182
rect 232 -186 235 -182
rect 249 -186 252 -182
rect 254 -186 264 -182
rect 266 -186 269 -182
rect 283 -186 286 -182
rect 288 -186 298 -182
rect 300 -186 303 -182
rect 317 -186 320 -182
rect 322 -186 332 -182
rect 334 -186 337 -182
rect 45 -262 48 -258
rect 50 -262 60 -258
rect 62 -262 65 -258
rect 79 -262 82 -258
rect 84 -262 94 -258
rect 96 -262 99 -258
rect 113 -262 116 -258
rect 118 -262 128 -258
rect 130 -262 133 -258
rect 147 -262 150 -258
rect 152 -262 162 -258
rect 164 -262 167 -258
rect 181 -262 184 -258
rect 186 -262 196 -258
rect 198 -262 201 -258
rect 215 -262 218 -258
rect 220 -262 230 -258
rect 232 -262 235 -258
rect 249 -262 252 -258
rect 254 -262 264 -258
rect 266 -262 269 -258
rect 283 -262 286 -258
rect 288 -262 298 -258
rect 300 -262 303 -258
rect 317 -262 320 -258
rect 322 -262 332 -258
rect 334 -262 337 -258
rect 45 -338 48 -334
rect 50 -338 60 -334
rect 62 -338 65 -334
rect 79 -338 82 -334
rect 84 -338 94 -334
rect 96 -338 99 -334
rect 113 -338 116 -334
rect 118 -338 128 -334
rect 130 -338 133 -334
rect 147 -338 150 -334
rect 152 -338 162 -334
rect 164 -338 167 -334
rect 181 -338 184 -334
rect 186 -338 196 -334
rect 198 -338 201 -334
rect 215 -338 218 -334
rect 220 -338 230 -334
rect 232 -338 235 -334
rect 249 -338 252 -334
rect 254 -338 264 -334
rect 266 -338 269 -334
rect 283 -338 286 -334
rect 288 -338 298 -334
rect 300 -338 303 -334
rect 317 -338 320 -334
rect 322 -338 332 -334
rect 334 -338 337 -334
rect 45 -414 48 -410
rect 50 -414 60 -410
rect 62 -414 65 -410
rect 79 -414 82 -410
rect 84 -414 94 -410
rect 96 -414 99 -410
rect 113 -414 116 -410
rect 118 -414 128 -410
rect 130 -414 133 -410
rect 147 -414 150 -410
rect 152 -414 162 -410
rect 164 -414 167 -410
rect 181 -414 184 -410
rect 186 -414 196 -410
rect 198 -414 201 -410
rect 215 -414 218 -410
rect 220 -414 230 -410
rect 232 -414 235 -410
rect 249 -414 252 -410
rect 254 -414 264 -410
rect 266 -414 269 -410
rect 283 -414 286 -410
rect 288 -414 298 -410
rect 300 -414 303 -410
rect 317 -414 320 -410
rect 322 -414 332 -410
rect 334 -414 337 -410
rect 45 -490 48 -486
rect 50 -490 60 -486
rect 62 -490 65 -486
rect 79 -490 82 -486
rect 84 -490 94 -486
rect 96 -490 99 -486
rect 113 -490 116 -486
rect 118 -490 128 -486
rect 130 -490 133 -486
rect 147 -490 150 -486
rect 152 -490 162 -486
rect 164 -490 167 -486
rect 181 -490 184 -486
rect 186 -490 196 -486
rect 198 -490 201 -486
rect 215 -490 218 -486
rect 220 -490 230 -486
rect 232 -490 235 -486
rect 249 -490 252 -486
rect 254 -490 264 -486
rect 266 -490 269 -486
rect 283 -490 286 -486
rect 288 -490 298 -486
rect 300 -490 303 -486
rect 317 -490 320 -486
rect 322 -490 332 -486
rect 334 -490 337 -486
rect 45 -566 48 -562
rect 50 -566 60 -562
rect 62 -566 65 -562
rect 79 -566 82 -562
rect 84 -566 94 -562
rect 96 -566 99 -562
rect 113 -566 116 -562
rect 118 -566 128 -562
rect 130 -566 133 -562
rect 147 -566 150 -562
rect 152 -566 162 -562
rect 164 -566 167 -562
rect 181 -566 184 -562
rect 186 -566 196 -562
rect 198 -566 201 -562
rect 215 -566 218 -562
rect 220 -566 230 -562
rect 232 -566 235 -562
rect 249 -566 252 -562
rect 254 -566 264 -562
rect 266 -566 269 -562
rect 283 -566 286 -562
rect 288 -566 298 -562
rect 300 -566 303 -562
rect 317 -566 320 -562
rect 322 -566 332 -562
rect 334 -566 337 -562
<< pdiffusion >>
rect 45 0 48 6
rect 50 0 53 6
rect 57 0 60 6
rect 62 0 65 6
rect 79 0 82 6
rect 84 0 87 6
rect 91 0 94 6
rect 96 0 99 6
rect 113 0 116 6
rect 118 0 121 6
rect 125 0 128 6
rect 130 0 133 6
rect 147 0 150 6
rect 152 0 155 6
rect 159 0 162 6
rect 164 0 167 6
rect 181 0 184 6
rect 186 0 189 6
rect 193 0 196 6
rect 198 0 201 6
rect 215 0 218 6
rect 220 0 223 6
rect 227 0 230 6
rect 232 0 235 6
rect 249 0 252 6
rect 254 0 257 6
rect 261 0 264 6
rect 266 0 269 6
rect 283 0 286 6
rect 288 0 291 6
rect 295 0 298 6
rect 300 0 303 6
rect 317 0 320 6
rect 322 0 325 6
rect 329 0 332 6
rect 334 0 337 6
rect 45 -76 48 -70
rect 50 -76 53 -70
rect 57 -76 60 -70
rect 62 -76 65 -70
rect 79 -76 82 -70
rect 84 -76 87 -70
rect 91 -76 94 -70
rect 96 -76 99 -70
rect 113 -76 116 -70
rect 118 -76 121 -70
rect 125 -76 128 -70
rect 130 -76 133 -70
rect 147 -76 150 -70
rect 152 -76 155 -70
rect 159 -76 162 -70
rect 164 -76 167 -70
rect 181 -76 184 -70
rect 186 -76 189 -70
rect 193 -76 196 -70
rect 198 -76 201 -70
rect 215 -76 218 -70
rect 220 -76 223 -70
rect 227 -76 230 -70
rect 232 -76 235 -70
rect 249 -76 252 -70
rect 254 -76 257 -70
rect 261 -76 264 -70
rect 266 -76 269 -70
rect 283 -76 286 -70
rect 288 -76 291 -70
rect 295 -76 298 -70
rect 300 -76 303 -70
rect 317 -76 320 -70
rect 322 -76 325 -70
rect 329 -76 332 -70
rect 334 -76 337 -70
rect 45 -152 48 -146
rect 50 -152 53 -146
rect 57 -152 60 -146
rect 62 -152 65 -146
rect 79 -152 82 -146
rect 84 -152 87 -146
rect 91 -152 94 -146
rect 96 -152 99 -146
rect 113 -152 116 -146
rect 118 -152 121 -146
rect 125 -152 128 -146
rect 130 -152 133 -146
rect 147 -152 150 -146
rect 152 -152 155 -146
rect 159 -152 162 -146
rect 164 -152 167 -146
rect 181 -152 184 -146
rect 186 -152 189 -146
rect 193 -152 196 -146
rect 198 -152 201 -146
rect 215 -152 218 -146
rect 220 -152 223 -146
rect 227 -152 230 -146
rect 232 -152 235 -146
rect 249 -152 252 -146
rect 254 -152 257 -146
rect 261 -152 264 -146
rect 266 -152 269 -146
rect 283 -152 286 -146
rect 288 -152 291 -146
rect 295 -152 298 -146
rect 300 -152 303 -146
rect 317 -152 320 -146
rect 322 -152 325 -146
rect 329 -152 332 -146
rect 334 -152 337 -146
rect 45 -228 48 -222
rect 50 -228 53 -222
rect 57 -228 60 -222
rect 62 -228 65 -222
rect 79 -228 82 -222
rect 84 -228 87 -222
rect 91 -228 94 -222
rect 96 -228 99 -222
rect 113 -228 116 -222
rect 118 -228 121 -222
rect 125 -228 128 -222
rect 130 -228 133 -222
rect 147 -228 150 -222
rect 152 -228 155 -222
rect 159 -228 162 -222
rect 164 -228 167 -222
rect 181 -228 184 -222
rect 186 -228 189 -222
rect 193 -228 196 -222
rect 198 -228 201 -222
rect 215 -228 218 -222
rect 220 -228 223 -222
rect 227 -228 230 -222
rect 232 -228 235 -222
rect 249 -228 252 -222
rect 254 -228 257 -222
rect 261 -228 264 -222
rect 266 -228 269 -222
rect 283 -228 286 -222
rect 288 -228 291 -222
rect 295 -228 298 -222
rect 300 -228 303 -222
rect 317 -228 320 -222
rect 322 -228 325 -222
rect 329 -228 332 -222
rect 334 -228 337 -222
rect 45 -304 48 -298
rect 50 -304 53 -298
rect 57 -304 60 -298
rect 62 -304 65 -298
rect 79 -304 82 -298
rect 84 -304 87 -298
rect 91 -304 94 -298
rect 96 -304 99 -298
rect 113 -304 116 -298
rect 118 -304 121 -298
rect 125 -304 128 -298
rect 130 -304 133 -298
rect 147 -304 150 -298
rect 152 -304 155 -298
rect 159 -304 162 -298
rect 164 -304 167 -298
rect 181 -304 184 -298
rect 186 -304 189 -298
rect 193 -304 196 -298
rect 198 -304 201 -298
rect 215 -304 218 -298
rect 220 -304 223 -298
rect 227 -304 230 -298
rect 232 -304 235 -298
rect 249 -304 252 -298
rect 254 -304 257 -298
rect 261 -304 264 -298
rect 266 -304 269 -298
rect 283 -304 286 -298
rect 288 -304 291 -298
rect 295 -304 298 -298
rect 300 -304 303 -298
rect 317 -304 320 -298
rect 322 -304 325 -298
rect 329 -304 332 -298
rect 334 -304 337 -298
rect 45 -380 48 -374
rect 50 -380 53 -374
rect 57 -380 60 -374
rect 62 -380 65 -374
rect 79 -380 82 -374
rect 84 -380 87 -374
rect 91 -380 94 -374
rect 96 -380 99 -374
rect 113 -380 116 -374
rect 118 -380 121 -374
rect 125 -380 128 -374
rect 130 -380 133 -374
rect 147 -380 150 -374
rect 152 -380 155 -374
rect 159 -380 162 -374
rect 164 -380 167 -374
rect 181 -380 184 -374
rect 186 -380 189 -374
rect 193 -380 196 -374
rect 198 -380 201 -374
rect 215 -380 218 -374
rect 220 -380 223 -374
rect 227 -380 230 -374
rect 232 -380 235 -374
rect 249 -380 252 -374
rect 254 -380 257 -374
rect 261 -380 264 -374
rect 266 -380 269 -374
rect 283 -380 286 -374
rect 288 -380 291 -374
rect 295 -380 298 -374
rect 300 -380 303 -374
rect 317 -380 320 -374
rect 322 -380 325 -374
rect 329 -380 332 -374
rect 334 -380 337 -374
rect 45 -456 48 -450
rect 50 -456 53 -450
rect 57 -456 60 -450
rect 62 -456 65 -450
rect 79 -456 82 -450
rect 84 -456 87 -450
rect 91 -456 94 -450
rect 96 -456 99 -450
rect 113 -456 116 -450
rect 118 -456 121 -450
rect 125 -456 128 -450
rect 130 -456 133 -450
rect 147 -456 150 -450
rect 152 -456 155 -450
rect 159 -456 162 -450
rect 164 -456 167 -450
rect 181 -456 184 -450
rect 186 -456 189 -450
rect 193 -456 196 -450
rect 198 -456 201 -450
rect 215 -456 218 -450
rect 220 -456 223 -450
rect 227 -456 230 -450
rect 232 -456 235 -450
rect 249 -456 252 -450
rect 254 -456 257 -450
rect 261 -456 264 -450
rect 266 -456 269 -450
rect 283 -456 286 -450
rect 288 -456 291 -450
rect 295 -456 298 -450
rect 300 -456 303 -450
rect 317 -456 320 -450
rect 322 -456 325 -450
rect 329 -456 332 -450
rect 334 -456 337 -450
rect 45 -532 48 -526
rect 50 -532 53 -526
rect 57 -532 60 -526
rect 62 -532 65 -526
rect 79 -532 82 -526
rect 84 -532 87 -526
rect 91 -532 94 -526
rect 96 -532 99 -526
rect 113 -532 116 -526
rect 118 -532 121 -526
rect 125 -532 128 -526
rect 130 -532 133 -526
rect 147 -532 150 -526
rect 152 -532 155 -526
rect 159 -532 162 -526
rect 164 -532 167 -526
rect 181 -532 184 -526
rect 186 -532 189 -526
rect 193 -532 196 -526
rect 198 -532 201 -526
rect 215 -532 218 -526
rect 220 -532 223 -526
rect 227 -532 230 -526
rect 232 -532 235 -526
rect 249 -532 252 -526
rect 254 -532 257 -526
rect 261 -532 264 -526
rect 266 -532 269 -526
rect 283 -532 286 -526
rect 288 -532 291 -526
rect 295 -532 298 -526
rect 300 -532 303 -526
rect 317 -532 320 -526
rect 322 -532 325 -526
rect 329 -532 332 -526
rect 334 -532 337 -526
<< ndcontact >>
rect 41 -34 45 -30
rect 65 -34 69 -30
rect 75 -34 79 -30
rect 99 -34 103 -30
rect 109 -34 113 -30
rect 133 -34 137 -30
rect 143 -34 147 -30
rect 167 -34 171 -30
rect 177 -34 181 -30
rect 201 -34 205 -30
rect 211 -34 215 -30
rect 235 -34 239 -30
rect 245 -34 249 -30
rect 269 -34 273 -30
rect 279 -34 283 -30
rect 303 -34 307 -30
rect 313 -34 317 -30
rect 337 -34 341 -30
rect 41 -110 45 -106
rect 65 -110 69 -106
rect 75 -110 79 -106
rect 99 -110 103 -106
rect 109 -110 113 -106
rect 133 -110 137 -106
rect 143 -110 147 -106
rect 167 -110 171 -106
rect 177 -110 181 -106
rect 201 -110 205 -106
rect 211 -110 215 -106
rect 235 -110 239 -106
rect 245 -110 249 -106
rect 269 -110 273 -106
rect 279 -110 283 -106
rect 303 -110 307 -106
rect 313 -110 317 -106
rect 337 -110 341 -106
rect 41 -186 45 -182
rect 65 -186 69 -182
rect 75 -186 79 -182
rect 99 -186 103 -182
rect 109 -186 113 -182
rect 133 -186 137 -182
rect 143 -186 147 -182
rect 167 -186 171 -182
rect 177 -186 181 -182
rect 201 -186 205 -182
rect 211 -186 215 -182
rect 235 -186 239 -182
rect 245 -186 249 -182
rect 269 -186 273 -182
rect 279 -186 283 -182
rect 303 -186 307 -182
rect 313 -186 317 -182
rect 337 -186 341 -182
rect 41 -262 45 -258
rect 65 -262 69 -258
rect 75 -262 79 -258
rect 99 -262 103 -258
rect 109 -262 113 -258
rect 133 -262 137 -258
rect 143 -262 147 -258
rect 167 -262 171 -258
rect 177 -262 181 -258
rect 201 -262 205 -258
rect 211 -262 215 -258
rect 235 -262 239 -258
rect 245 -262 249 -258
rect 269 -262 273 -258
rect 279 -262 283 -258
rect 303 -262 307 -258
rect 313 -262 317 -258
rect 337 -262 341 -258
rect 41 -338 45 -334
rect 65 -338 69 -334
rect 75 -338 79 -334
rect 99 -338 103 -334
rect 109 -338 113 -334
rect 133 -338 137 -334
rect 143 -338 147 -334
rect 167 -338 171 -334
rect 177 -338 181 -334
rect 201 -338 205 -334
rect 211 -338 215 -334
rect 235 -338 239 -334
rect 245 -338 249 -334
rect 269 -338 273 -334
rect 279 -338 283 -334
rect 303 -338 307 -334
rect 313 -338 317 -334
rect 337 -338 341 -334
rect 41 -414 45 -410
rect 65 -414 69 -410
rect 75 -414 79 -410
rect 99 -414 103 -410
rect 109 -414 113 -410
rect 133 -414 137 -410
rect 143 -414 147 -410
rect 167 -414 171 -410
rect 177 -414 181 -410
rect 201 -414 205 -410
rect 211 -414 215 -410
rect 235 -414 239 -410
rect 245 -414 249 -410
rect 269 -414 273 -410
rect 279 -414 283 -410
rect 303 -414 307 -410
rect 313 -414 317 -410
rect 337 -414 341 -410
rect 41 -490 45 -486
rect 65 -490 69 -486
rect 75 -490 79 -486
rect 99 -490 103 -486
rect 109 -490 113 -486
rect 133 -490 137 -486
rect 143 -490 147 -486
rect 167 -490 171 -486
rect 177 -490 181 -486
rect 201 -490 205 -486
rect 211 -490 215 -486
rect 235 -490 239 -486
rect 245 -490 249 -486
rect 269 -490 273 -486
rect 279 -490 283 -486
rect 303 -490 307 -486
rect 313 -490 317 -486
rect 337 -490 341 -486
rect 41 -566 45 -562
rect 65 -566 69 -562
rect 75 -566 79 -562
rect 99 -566 103 -562
rect 109 -566 113 -562
rect 133 -566 137 -562
rect 143 -566 147 -562
rect 167 -566 171 -562
rect 177 -566 181 -562
rect 201 -566 205 -562
rect 211 -566 215 -562
rect 235 -566 239 -562
rect 245 -566 249 -562
rect 269 -566 273 -562
rect 279 -566 283 -562
rect 303 -566 307 -562
rect 313 -566 317 -562
rect 337 -566 341 -562
<< pdcontact >>
rect 41 0 45 6
rect 53 0 57 6
rect 65 0 69 6
rect 75 0 79 6
rect 87 0 91 6
rect 99 0 103 6
rect 109 0 113 6
rect 121 0 125 6
rect 133 0 137 6
rect 143 0 147 6
rect 155 0 159 6
rect 167 0 171 6
rect 177 0 181 6
rect 189 0 193 6
rect 201 0 205 6
rect 211 0 215 6
rect 223 0 227 6
rect 235 0 239 6
rect 245 0 249 6
rect 257 0 261 6
rect 269 0 273 6
rect 279 0 283 6
rect 291 0 295 6
rect 303 0 307 6
rect 313 0 317 6
rect 325 0 329 6
rect 337 0 341 6
rect 41 -76 45 -70
rect 53 -76 57 -70
rect 65 -76 69 -70
rect 75 -76 79 -70
rect 87 -76 91 -70
rect 99 -76 103 -70
rect 109 -76 113 -70
rect 121 -76 125 -70
rect 133 -76 137 -70
rect 143 -76 147 -70
rect 155 -76 159 -70
rect 167 -76 171 -70
rect 177 -76 181 -70
rect 189 -76 193 -70
rect 201 -76 205 -70
rect 211 -76 215 -70
rect 223 -76 227 -70
rect 235 -76 239 -70
rect 245 -76 249 -70
rect 257 -76 261 -70
rect 269 -76 273 -70
rect 279 -76 283 -70
rect 291 -76 295 -70
rect 303 -76 307 -70
rect 313 -76 317 -70
rect 325 -76 329 -70
rect 337 -76 341 -70
rect 41 -152 45 -146
rect 53 -152 57 -146
rect 65 -152 69 -146
rect 75 -152 79 -146
rect 87 -152 91 -146
rect 99 -152 103 -146
rect 109 -152 113 -146
rect 121 -152 125 -146
rect 133 -152 137 -146
rect 143 -152 147 -146
rect 155 -152 159 -146
rect 167 -152 171 -146
rect 177 -152 181 -146
rect 189 -152 193 -146
rect 201 -152 205 -146
rect 211 -152 215 -146
rect 223 -152 227 -146
rect 235 -152 239 -146
rect 245 -152 249 -146
rect 257 -152 261 -146
rect 269 -152 273 -146
rect 279 -152 283 -146
rect 291 -152 295 -146
rect 303 -152 307 -146
rect 313 -152 317 -146
rect 325 -152 329 -146
rect 337 -152 341 -146
rect 41 -228 45 -222
rect 53 -228 57 -222
rect 65 -228 69 -222
rect 75 -228 79 -222
rect 87 -228 91 -222
rect 99 -228 103 -222
rect 109 -228 113 -222
rect 121 -228 125 -222
rect 133 -228 137 -222
rect 143 -228 147 -222
rect 155 -228 159 -222
rect 167 -228 171 -222
rect 177 -228 181 -222
rect 189 -228 193 -222
rect 201 -228 205 -222
rect 211 -228 215 -222
rect 223 -228 227 -222
rect 235 -228 239 -222
rect 245 -228 249 -222
rect 257 -228 261 -222
rect 269 -228 273 -222
rect 279 -228 283 -222
rect 291 -228 295 -222
rect 303 -228 307 -222
rect 313 -228 317 -222
rect 325 -228 329 -222
rect 337 -228 341 -222
rect 41 -304 45 -298
rect 53 -304 57 -298
rect 65 -304 69 -298
rect 75 -304 79 -298
rect 87 -304 91 -298
rect 99 -304 103 -298
rect 109 -304 113 -298
rect 121 -304 125 -298
rect 133 -304 137 -298
rect 143 -304 147 -298
rect 155 -304 159 -298
rect 167 -304 171 -298
rect 177 -304 181 -298
rect 189 -304 193 -298
rect 201 -304 205 -298
rect 211 -304 215 -298
rect 223 -304 227 -298
rect 235 -304 239 -298
rect 245 -304 249 -298
rect 257 -304 261 -298
rect 269 -304 273 -298
rect 279 -304 283 -298
rect 291 -304 295 -298
rect 303 -304 307 -298
rect 313 -304 317 -298
rect 325 -304 329 -298
rect 337 -304 341 -298
rect 41 -380 45 -374
rect 53 -380 57 -374
rect 65 -380 69 -374
rect 75 -380 79 -374
rect 87 -380 91 -374
rect 99 -380 103 -374
rect 109 -380 113 -374
rect 121 -380 125 -374
rect 133 -380 137 -374
rect 143 -380 147 -374
rect 155 -380 159 -374
rect 167 -380 171 -374
rect 177 -380 181 -374
rect 189 -380 193 -374
rect 201 -380 205 -374
rect 211 -380 215 -374
rect 223 -380 227 -374
rect 235 -380 239 -374
rect 245 -380 249 -374
rect 257 -380 261 -374
rect 269 -380 273 -374
rect 279 -380 283 -374
rect 291 -380 295 -374
rect 303 -380 307 -374
rect 313 -380 317 -374
rect 325 -380 329 -374
rect 337 -380 341 -374
rect 41 -456 45 -450
rect 53 -456 57 -450
rect 65 -456 69 -450
rect 75 -456 79 -450
rect 87 -456 91 -450
rect 99 -456 103 -450
rect 109 -456 113 -450
rect 121 -456 125 -450
rect 133 -456 137 -450
rect 143 -456 147 -450
rect 155 -456 159 -450
rect 167 -456 171 -450
rect 177 -456 181 -450
rect 189 -456 193 -450
rect 201 -456 205 -450
rect 211 -456 215 -450
rect 223 -456 227 -450
rect 235 -456 239 -450
rect 245 -456 249 -450
rect 257 -456 261 -450
rect 269 -456 273 -450
rect 279 -456 283 -450
rect 291 -456 295 -450
rect 303 -456 307 -450
rect 313 -456 317 -450
rect 325 -456 329 -450
rect 337 -456 341 -450
rect 41 -532 45 -526
rect 53 -532 57 -526
rect 65 -532 69 -526
rect 75 -532 79 -526
rect 87 -532 91 -526
rect 99 -532 103 -526
rect 109 -532 113 -526
rect 121 -532 125 -526
rect 133 -532 137 -526
rect 143 -532 147 -526
rect 155 -532 159 -526
rect 167 -532 171 -526
rect 177 -532 181 -526
rect 189 -532 193 -526
rect 201 -532 205 -526
rect 211 -532 215 -526
rect 223 -532 227 -526
rect 235 -532 239 -526
rect 245 -532 249 -526
rect 257 -532 261 -526
rect 269 -532 273 -526
rect 279 -532 283 -526
rect 291 -532 295 -526
rect 303 -532 307 -526
rect 313 -532 317 -526
rect 325 -532 329 -526
rect 337 -532 341 -526
<< polysilicon >>
rect 48 6 50 9
rect 60 6 62 9
rect 82 6 84 9
rect 94 6 96 9
rect 116 6 118 9
rect 128 6 130 9
rect 150 6 152 9
rect 162 6 164 9
rect 184 6 186 9
rect 196 6 198 9
rect 218 6 220 9
rect 230 6 232 9
rect 252 6 254 9
rect 264 6 266 9
rect 286 6 288 9
rect 298 6 300 9
rect 320 6 322 9
rect 332 6 334 9
rect 48 -30 50 0
rect 60 -30 62 0
rect 82 -30 84 0
rect 94 -30 96 0
rect 116 -30 118 0
rect 128 -30 130 0
rect 150 -30 152 0
rect 162 -30 164 0
rect 184 -30 186 0
rect 196 -30 198 0
rect 218 -30 220 0
rect 230 -30 232 0
rect 252 -30 254 0
rect 264 -30 266 0
rect 286 -30 288 0
rect 298 -30 300 0
rect 320 -30 322 0
rect 332 -30 334 0
rect 48 -37 50 -34
rect 60 -37 62 -34
rect 82 -37 84 -34
rect 94 -38 96 -34
rect 116 -37 118 -34
rect 128 -37 130 -34
rect 150 -37 152 -34
rect 162 -37 164 -34
rect 184 -37 186 -34
rect 196 -37 198 -34
rect 218 -37 220 -34
rect 230 -37 232 -34
rect 252 -37 254 -34
rect 264 -37 266 -34
rect 286 -37 288 -34
rect 298 -37 300 -34
rect 320 -37 322 -34
rect 332 -37 334 -34
rect 48 -70 50 -67
rect 60 -70 62 -67
rect 82 -70 84 -67
rect 94 -70 96 -67
rect 116 -70 118 -67
rect 128 -70 130 -67
rect 150 -70 152 -67
rect 162 -70 164 -67
rect 184 -70 186 -67
rect 196 -70 198 -67
rect 218 -70 220 -67
rect 230 -70 232 -67
rect 252 -70 254 -67
rect 264 -70 266 -67
rect 286 -70 288 -67
rect 298 -70 300 -67
rect 320 -70 322 -67
rect 332 -70 334 -67
rect 48 -106 50 -76
rect 60 -106 62 -76
rect 82 -106 84 -76
rect 94 -106 96 -76
rect 116 -106 118 -76
rect 128 -106 130 -76
rect 150 -106 152 -76
rect 162 -106 164 -76
rect 184 -106 186 -76
rect 196 -106 198 -76
rect 218 -106 220 -76
rect 230 -106 232 -76
rect 252 -106 254 -76
rect 264 -106 266 -76
rect 286 -106 288 -76
rect 298 -106 300 -76
rect 320 -106 322 -76
rect 332 -106 334 -76
rect 48 -113 50 -110
rect 60 -113 62 -110
rect 82 -113 84 -110
rect 94 -114 96 -110
rect 116 -113 118 -110
rect 128 -113 130 -110
rect 150 -113 152 -110
rect 162 -113 164 -110
rect 184 -113 186 -110
rect 196 -113 198 -110
rect 218 -113 220 -110
rect 230 -113 232 -110
rect 252 -113 254 -110
rect 264 -113 266 -110
rect 286 -113 288 -110
rect 298 -113 300 -110
rect 320 -113 322 -110
rect 332 -113 334 -110
rect 48 -146 50 -143
rect 60 -146 62 -143
rect 82 -146 84 -143
rect 94 -146 96 -143
rect 116 -146 118 -143
rect 128 -146 130 -143
rect 150 -146 152 -143
rect 162 -146 164 -143
rect 184 -146 186 -143
rect 196 -146 198 -143
rect 218 -146 220 -143
rect 230 -146 232 -143
rect 252 -146 254 -143
rect 264 -146 266 -143
rect 286 -146 288 -143
rect 298 -146 300 -143
rect 320 -146 322 -143
rect 332 -146 334 -143
rect 48 -182 50 -152
rect 60 -182 62 -152
rect 82 -182 84 -152
rect 94 -182 96 -152
rect 116 -182 118 -152
rect 128 -182 130 -152
rect 150 -182 152 -152
rect 162 -182 164 -152
rect 184 -182 186 -152
rect 196 -182 198 -152
rect 218 -182 220 -152
rect 230 -182 232 -152
rect 252 -182 254 -152
rect 264 -182 266 -152
rect 286 -182 288 -152
rect 298 -182 300 -152
rect 320 -182 322 -152
rect 332 -182 334 -152
rect 48 -189 50 -186
rect 60 -189 62 -186
rect 82 -189 84 -186
rect 94 -190 96 -186
rect 116 -189 118 -186
rect 128 -189 130 -186
rect 150 -189 152 -186
rect 162 -189 164 -186
rect 184 -189 186 -186
rect 196 -189 198 -186
rect 218 -189 220 -186
rect 230 -189 232 -186
rect 252 -189 254 -186
rect 264 -189 266 -186
rect 286 -189 288 -186
rect 298 -189 300 -186
rect 320 -189 322 -186
rect 332 -189 334 -186
rect 48 -222 50 -219
rect 60 -222 62 -219
rect 82 -222 84 -219
rect 94 -222 96 -219
rect 116 -222 118 -219
rect 128 -222 130 -219
rect 150 -222 152 -219
rect 162 -222 164 -219
rect 184 -222 186 -219
rect 196 -222 198 -219
rect 218 -222 220 -219
rect 230 -222 232 -219
rect 252 -222 254 -219
rect 264 -222 266 -219
rect 286 -222 288 -219
rect 298 -222 300 -219
rect 320 -222 322 -219
rect 332 -222 334 -219
rect 48 -258 50 -228
rect 60 -258 62 -228
rect 82 -258 84 -228
rect 94 -258 96 -228
rect 116 -258 118 -228
rect 128 -258 130 -228
rect 150 -258 152 -228
rect 162 -258 164 -228
rect 184 -258 186 -228
rect 196 -258 198 -228
rect 218 -258 220 -228
rect 230 -258 232 -228
rect 252 -258 254 -228
rect 264 -258 266 -228
rect 286 -258 288 -228
rect 298 -258 300 -228
rect 320 -258 322 -228
rect 332 -258 334 -228
rect 48 -265 50 -262
rect 60 -265 62 -262
rect 82 -265 84 -262
rect 94 -266 96 -262
rect 116 -265 118 -262
rect 128 -265 130 -262
rect 150 -265 152 -262
rect 162 -265 164 -262
rect 184 -265 186 -262
rect 196 -265 198 -262
rect 218 -265 220 -262
rect 230 -265 232 -262
rect 252 -265 254 -262
rect 264 -265 266 -262
rect 286 -265 288 -262
rect 298 -265 300 -262
rect 320 -265 322 -262
rect 332 -265 334 -262
rect 48 -298 50 -295
rect 60 -298 62 -295
rect 82 -298 84 -295
rect 94 -298 96 -295
rect 116 -298 118 -295
rect 128 -298 130 -295
rect 150 -298 152 -295
rect 162 -298 164 -295
rect 184 -298 186 -295
rect 196 -298 198 -295
rect 218 -298 220 -295
rect 230 -298 232 -295
rect 252 -298 254 -295
rect 264 -298 266 -295
rect 286 -298 288 -295
rect 298 -298 300 -295
rect 320 -298 322 -295
rect 332 -298 334 -295
rect 48 -334 50 -304
rect 60 -334 62 -304
rect 82 -334 84 -304
rect 94 -334 96 -304
rect 116 -334 118 -304
rect 128 -334 130 -304
rect 150 -334 152 -304
rect 162 -334 164 -304
rect 184 -334 186 -304
rect 196 -334 198 -304
rect 218 -334 220 -304
rect 230 -334 232 -304
rect 252 -334 254 -304
rect 264 -334 266 -304
rect 286 -334 288 -304
rect 298 -334 300 -304
rect 320 -334 322 -304
rect 332 -334 334 -304
rect 48 -341 50 -338
rect 60 -341 62 -338
rect 82 -341 84 -338
rect 94 -342 96 -338
rect 116 -341 118 -338
rect 128 -341 130 -338
rect 150 -341 152 -338
rect 162 -341 164 -338
rect 184 -341 186 -338
rect 196 -341 198 -338
rect 218 -341 220 -338
rect 230 -341 232 -338
rect 252 -341 254 -338
rect 264 -341 266 -338
rect 286 -341 288 -338
rect 298 -341 300 -338
rect 320 -341 322 -338
rect 332 -341 334 -338
rect 48 -374 50 -371
rect 60 -374 62 -371
rect 82 -374 84 -371
rect 94 -374 96 -371
rect 116 -374 118 -371
rect 128 -374 130 -371
rect 150 -374 152 -371
rect 162 -374 164 -371
rect 184 -374 186 -371
rect 196 -374 198 -371
rect 218 -374 220 -371
rect 230 -374 232 -371
rect 252 -374 254 -371
rect 264 -374 266 -371
rect 286 -374 288 -371
rect 298 -374 300 -371
rect 320 -374 322 -371
rect 332 -374 334 -371
rect 48 -410 50 -380
rect 60 -410 62 -380
rect 82 -410 84 -380
rect 94 -410 96 -380
rect 116 -410 118 -380
rect 128 -410 130 -380
rect 150 -410 152 -380
rect 162 -410 164 -380
rect 184 -410 186 -380
rect 196 -410 198 -380
rect 218 -410 220 -380
rect 230 -410 232 -380
rect 252 -410 254 -380
rect 264 -410 266 -380
rect 286 -410 288 -380
rect 298 -410 300 -380
rect 320 -410 322 -380
rect 332 -410 334 -380
rect 48 -417 50 -414
rect 60 -417 62 -414
rect 82 -417 84 -414
rect 94 -418 96 -414
rect 116 -417 118 -414
rect 128 -417 130 -414
rect 150 -417 152 -414
rect 162 -417 164 -414
rect 184 -417 186 -414
rect 196 -417 198 -414
rect 218 -417 220 -414
rect 230 -417 232 -414
rect 252 -417 254 -414
rect 264 -417 266 -414
rect 286 -417 288 -414
rect 298 -417 300 -414
rect 320 -417 322 -414
rect 332 -417 334 -414
rect 48 -450 50 -447
rect 60 -450 62 -447
rect 82 -450 84 -447
rect 94 -450 96 -447
rect 116 -450 118 -447
rect 128 -450 130 -447
rect 150 -450 152 -447
rect 162 -450 164 -447
rect 184 -450 186 -447
rect 196 -450 198 -447
rect 218 -450 220 -447
rect 230 -450 232 -447
rect 252 -450 254 -447
rect 264 -450 266 -447
rect 286 -450 288 -447
rect 298 -450 300 -447
rect 320 -450 322 -447
rect 332 -450 334 -447
rect 48 -486 50 -456
rect 60 -486 62 -456
rect 82 -486 84 -456
rect 94 -486 96 -456
rect 116 -486 118 -456
rect 128 -486 130 -456
rect 150 -486 152 -456
rect 162 -486 164 -456
rect 184 -486 186 -456
rect 196 -486 198 -456
rect 218 -486 220 -456
rect 230 -486 232 -456
rect 252 -486 254 -456
rect 264 -486 266 -456
rect 286 -486 288 -456
rect 298 -486 300 -456
rect 320 -486 322 -456
rect 332 -486 334 -456
rect 48 -493 50 -490
rect 60 -493 62 -490
rect 82 -493 84 -490
rect 94 -494 96 -490
rect 116 -493 118 -490
rect 128 -493 130 -490
rect 150 -493 152 -490
rect 162 -493 164 -490
rect 184 -493 186 -490
rect 196 -493 198 -490
rect 218 -493 220 -490
rect 230 -493 232 -490
rect 252 -493 254 -490
rect 264 -493 266 -490
rect 286 -493 288 -490
rect 298 -493 300 -490
rect 320 -493 322 -490
rect 332 -493 334 -490
rect 48 -526 50 -523
rect 60 -526 62 -523
rect 82 -526 84 -523
rect 94 -526 96 -523
rect 116 -526 118 -523
rect 128 -526 130 -523
rect 150 -526 152 -523
rect 162 -526 164 -523
rect 184 -526 186 -523
rect 196 -526 198 -523
rect 218 -526 220 -523
rect 230 -526 232 -523
rect 252 -526 254 -523
rect 264 -526 266 -523
rect 286 -526 288 -523
rect 298 -526 300 -523
rect 320 -526 322 -523
rect 332 -526 334 -523
rect 48 -562 50 -532
rect 60 -562 62 -532
rect 82 -562 84 -532
rect 94 -562 96 -532
rect 116 -562 118 -532
rect 128 -562 130 -532
rect 150 -562 152 -532
rect 162 -562 164 -532
rect 184 -562 186 -532
rect 196 -562 198 -532
rect 218 -562 220 -532
rect 230 -562 232 -532
rect 252 -562 254 -532
rect 264 -562 266 -532
rect 286 -562 288 -532
rect 298 -562 300 -532
rect 320 -562 322 -532
rect 332 -562 334 -532
rect 48 -569 50 -566
rect 60 -569 62 -566
rect 82 -569 84 -566
rect 94 -570 96 -566
rect 116 -569 118 -566
rect 128 -569 130 -566
rect 150 -569 152 -566
rect 162 -569 164 -566
rect 184 -569 186 -566
rect 196 -569 198 -566
rect 218 -569 220 -566
rect 230 -569 232 -566
rect 252 -569 254 -566
rect 264 -569 266 -566
rect 286 -569 288 -566
rect 298 -569 300 -566
rect 320 -569 322 -566
rect 332 -569 334 -566
<< polycontact >>
rect 44 -21 48 -17
rect 56 -21 60 -17
rect 78 -14 82 -10
rect 90 -28 94 -24
rect 124 -14 128 -10
rect 146 -26 150 -22
rect 158 -21 162 -17
rect 180 -14 184 -10
rect 192 -26 196 -22
rect 214 -17 218 -13
rect 226 -27 230 -23
rect 248 -8 252 -4
rect 260 -28 264 -24
rect 282 -10 286 -6
rect 294 -25 298 -21
rect 316 -16 320 -12
rect 116 -41 120 -37
rect 332 -41 336 -37
rect 44 -97 48 -93
rect 56 -97 60 -93
rect 78 -90 82 -86
rect 90 -104 94 -100
rect 124 -90 128 -86
rect 146 -102 150 -98
rect 158 -97 162 -93
rect 180 -90 184 -86
rect 192 -102 196 -98
rect 214 -93 218 -89
rect 226 -103 230 -99
rect 248 -84 252 -80
rect 260 -104 264 -100
rect 282 -86 286 -82
rect 294 -101 298 -97
rect 316 -92 320 -88
rect 116 -117 120 -113
rect 332 -117 336 -113
rect 44 -173 48 -169
rect 56 -173 60 -169
rect 78 -166 82 -162
rect 90 -180 94 -176
rect 124 -166 128 -162
rect 146 -178 150 -174
rect 158 -173 162 -169
rect 180 -166 184 -162
rect 192 -178 196 -174
rect 214 -169 218 -165
rect 226 -179 230 -175
rect 248 -160 252 -156
rect 260 -180 264 -176
rect 282 -162 286 -158
rect 294 -177 298 -173
rect 316 -168 320 -164
rect 116 -193 120 -189
rect 332 -193 336 -189
rect 44 -249 48 -245
rect 56 -249 60 -245
rect 78 -242 82 -238
rect 90 -256 94 -252
rect 124 -242 128 -238
rect 146 -254 150 -250
rect 158 -249 162 -245
rect 180 -242 184 -238
rect 192 -254 196 -250
rect 214 -245 218 -241
rect 226 -255 230 -251
rect 248 -236 252 -232
rect 260 -256 264 -252
rect 282 -238 286 -234
rect 294 -253 298 -249
rect 316 -244 320 -240
rect 116 -269 120 -265
rect 332 -269 336 -265
rect 44 -325 48 -321
rect 56 -325 60 -321
rect 78 -318 82 -314
rect 90 -332 94 -328
rect 124 -318 128 -314
rect 146 -330 150 -326
rect 158 -325 162 -321
rect 180 -318 184 -314
rect 192 -330 196 -326
rect 214 -321 218 -317
rect 226 -331 230 -327
rect 248 -312 252 -308
rect 260 -332 264 -328
rect 282 -314 286 -310
rect 294 -329 298 -325
rect 316 -320 320 -316
rect 116 -345 120 -341
rect 332 -345 336 -341
rect 44 -401 48 -397
rect 56 -401 60 -397
rect 78 -394 82 -390
rect 90 -408 94 -404
rect 124 -394 128 -390
rect 146 -406 150 -402
rect 158 -401 162 -397
rect 180 -394 184 -390
rect 192 -406 196 -402
rect 214 -397 218 -393
rect 226 -407 230 -403
rect 248 -388 252 -384
rect 260 -408 264 -404
rect 282 -390 286 -386
rect 294 -405 298 -401
rect 316 -396 320 -392
rect 116 -421 120 -417
rect 332 -421 336 -417
rect 44 -477 48 -473
rect 56 -477 60 -473
rect 78 -470 82 -466
rect 90 -484 94 -480
rect 124 -470 128 -466
rect 146 -482 150 -478
rect 158 -477 162 -473
rect 180 -470 184 -466
rect 192 -482 196 -478
rect 214 -473 218 -469
rect 226 -483 230 -479
rect 248 -464 252 -460
rect 260 -484 264 -480
rect 282 -466 286 -462
rect 294 -481 298 -477
rect 316 -472 320 -468
rect 116 -497 120 -493
rect 332 -497 336 -493
rect 44 -553 48 -549
rect 56 -553 60 -549
rect 78 -546 82 -542
rect 90 -560 94 -556
rect 124 -546 128 -542
rect 146 -558 150 -554
rect 158 -553 162 -549
rect 180 -546 184 -542
rect 192 -558 196 -554
rect 214 -549 218 -545
rect 226 -559 230 -555
rect 248 -540 252 -536
rect 260 -560 264 -556
rect 282 -542 286 -538
rect 294 -557 298 -553
rect 316 -548 320 -544
rect 116 -573 120 -569
rect 332 -573 336 -569
<< metal1 >>
rect -14 -577 -6 27
rect 2 25 10 27
rect 2 16 347 25
rect 2 -54 10 16
rect 28 4 35 8
rect 41 6 45 16
rect 65 6 69 16
rect 75 6 79 16
rect 99 6 103 16
rect 109 6 113 16
rect 133 6 137 16
rect 143 6 147 16
rect 167 6 171 16
rect 177 6 181 16
rect 201 6 205 16
rect 211 6 215 16
rect 235 6 239 16
rect 245 6 249 16
rect 269 6 273 16
rect 279 6 283 16
rect 303 6 307 16
rect 313 6 317 16
rect 337 6 341 16
rect 28 -13 35 -9
rect 53 -10 57 0
rect 53 -14 65 -10
rect 70 -14 78 -10
rect 87 -11 91 0
rect 121 -3 125 0
rect 121 -7 137 -3
rect 28 -21 35 -17
rect 40 -21 44 -17
rect 65 -30 69 -14
rect 87 -15 103 -11
rect 99 -30 103 -15
rect 133 -30 137 -7
rect 155 -10 159 0
rect 155 -14 171 -10
rect 176 -14 180 -10
rect 189 -13 193 0
rect 223 -12 227 0
rect 257 -6 261 0
rect 291 -4 295 0
rect 257 -10 282 -6
rect 291 -8 315 -4
rect 167 -30 171 -14
rect 189 -17 205 -13
rect 210 -17 214 -13
rect 223 -16 244 -12
rect 201 -30 205 -17
rect 213 -27 226 -23
rect 235 -30 239 -16
rect 269 -30 273 -10
rect 284 -25 294 -21
rect 303 -30 307 -8
rect 325 -12 329 0
rect 311 -16 316 -12
rect 325 -16 342 -12
rect 311 -19 315 -16
rect 337 -30 341 -16
rect 41 -45 45 -34
rect 75 -45 79 -34
rect 109 -45 113 -34
rect 143 -45 147 -34
rect 177 -45 181 -34
rect 211 -45 215 -34
rect 245 -45 249 -34
rect 279 -45 283 -34
rect 313 -45 317 -34
rect 329 -41 332 -37
rect 24 -46 346 -45
rect 24 -50 347 -46
rect 24 -51 346 -50
rect 2 -62 347 -54
rect 2 -131 10 -62
rect 41 -70 45 -62
rect 65 -70 69 -62
rect 75 -70 79 -62
rect 99 -70 103 -62
rect 109 -70 113 -62
rect 133 -70 137 -62
rect 143 -70 147 -62
rect 167 -70 171 -62
rect 177 -70 181 -62
rect 201 -70 205 -62
rect 211 -70 215 -62
rect 235 -70 239 -62
rect 245 -70 249 -62
rect 269 -70 273 -62
rect 279 -70 283 -62
rect 303 -70 307 -62
rect 313 -70 317 -62
rect 337 -70 341 -62
rect 28 -89 35 -85
rect 53 -86 57 -76
rect 53 -90 65 -86
rect 70 -90 78 -86
rect 87 -87 91 -76
rect 121 -79 125 -76
rect 121 -83 137 -79
rect 28 -97 35 -93
rect 40 -97 44 -93
rect 65 -106 69 -90
rect 87 -91 103 -87
rect 99 -106 103 -91
rect 133 -106 137 -83
rect 155 -86 159 -76
rect 155 -90 171 -86
rect 176 -90 180 -86
rect 189 -89 193 -76
rect 223 -88 227 -76
rect 257 -82 261 -76
rect 291 -80 295 -76
rect 257 -86 282 -82
rect 291 -84 315 -80
rect 167 -106 171 -90
rect 189 -93 205 -89
rect 210 -93 214 -89
rect 223 -92 244 -88
rect 201 -106 205 -93
rect 213 -103 226 -99
rect 235 -106 239 -92
rect 269 -106 273 -86
rect 284 -101 294 -97
rect 303 -106 307 -84
rect 325 -88 329 -76
rect 311 -92 316 -88
rect 325 -92 342 -88
rect 311 -95 315 -92
rect 337 -106 341 -92
rect 41 -121 45 -110
rect 75 -121 79 -110
rect 109 -121 113 -110
rect 143 -121 147 -110
rect 177 -121 181 -110
rect 211 -121 215 -110
rect 245 -121 249 -110
rect 279 -121 283 -110
rect 313 -121 317 -110
rect 329 -117 332 -113
rect 24 -128 347 -121
rect 2 -139 347 -131
rect 2 -207 10 -139
rect 30 -140 35 -139
rect 41 -146 45 -139
rect 65 -146 69 -139
rect 75 -146 79 -139
rect 99 -146 103 -139
rect 109 -146 113 -139
rect 133 -146 137 -139
rect 143 -146 147 -139
rect 167 -146 171 -139
rect 177 -146 181 -139
rect 201 -146 205 -139
rect 211 -146 215 -139
rect 235 -146 239 -139
rect 245 -146 249 -139
rect 269 -146 273 -139
rect 279 -146 283 -139
rect 303 -146 307 -139
rect 313 -146 317 -139
rect 337 -146 341 -139
rect 28 -165 35 -161
rect 53 -162 57 -152
rect 53 -166 65 -162
rect 70 -166 78 -162
rect 87 -163 91 -152
rect 121 -155 125 -152
rect 121 -159 137 -155
rect 28 -173 35 -169
rect 40 -173 44 -169
rect 65 -182 69 -166
rect 87 -167 103 -163
rect 99 -182 103 -167
rect 133 -182 137 -159
rect 155 -162 159 -152
rect 155 -166 171 -162
rect 176 -166 180 -162
rect 189 -165 193 -152
rect 223 -164 227 -152
rect 257 -158 261 -152
rect 291 -156 295 -152
rect 257 -162 282 -158
rect 291 -160 315 -156
rect 167 -182 171 -166
rect 189 -169 205 -165
rect 210 -169 214 -165
rect 223 -168 244 -164
rect 201 -182 205 -169
rect 213 -179 226 -175
rect 235 -182 239 -168
rect 269 -182 273 -162
rect 284 -177 294 -173
rect 303 -182 307 -160
rect 325 -164 329 -152
rect 311 -168 316 -164
rect 325 -168 342 -164
rect 311 -171 315 -168
rect 337 -182 341 -168
rect 41 -197 45 -186
rect 75 -197 79 -186
rect 109 -197 113 -186
rect 143 -197 147 -186
rect 177 -197 181 -186
rect 211 -197 215 -186
rect 245 -197 249 -186
rect 279 -197 283 -186
rect 313 -197 317 -186
rect 329 -193 332 -189
rect 24 -204 347 -197
rect 2 -215 347 -207
rect 2 -284 10 -215
rect 30 -220 35 -215
rect 41 -222 45 -215
rect 65 -222 69 -215
rect 75 -222 79 -215
rect 99 -222 103 -215
rect 109 -222 113 -215
rect 133 -222 137 -215
rect 143 -222 147 -215
rect 167 -222 171 -215
rect 177 -222 181 -215
rect 201 -222 205 -215
rect 211 -222 215 -215
rect 235 -222 239 -215
rect 245 -222 249 -215
rect 269 -222 273 -215
rect 279 -222 283 -215
rect 303 -222 307 -215
rect 313 -222 317 -215
rect 337 -222 341 -215
rect 28 -241 35 -237
rect 53 -238 57 -228
rect 53 -242 65 -238
rect 70 -242 78 -238
rect 87 -239 91 -228
rect 121 -231 125 -228
rect 121 -235 137 -231
rect 28 -249 35 -245
rect 40 -249 44 -245
rect 65 -258 69 -242
rect 87 -243 103 -239
rect 99 -258 103 -243
rect 133 -258 137 -235
rect 155 -238 159 -228
rect 155 -242 171 -238
rect 176 -242 180 -238
rect 189 -241 193 -228
rect 223 -240 227 -228
rect 257 -234 261 -228
rect 291 -232 295 -228
rect 257 -238 282 -234
rect 291 -236 315 -232
rect 167 -258 171 -242
rect 189 -245 205 -241
rect 210 -245 214 -241
rect 223 -244 244 -240
rect 201 -258 205 -245
rect 213 -255 226 -251
rect 235 -258 239 -244
rect 269 -258 273 -238
rect 284 -253 294 -249
rect 303 -258 307 -236
rect 325 -240 329 -228
rect 311 -244 316 -240
rect 325 -244 342 -240
rect 311 -247 315 -244
rect 337 -258 341 -244
rect 41 -273 45 -262
rect 75 -273 79 -262
rect 109 -273 113 -262
rect 143 -273 147 -262
rect 177 -273 181 -262
rect 211 -273 215 -262
rect 245 -273 249 -262
rect 279 -273 283 -262
rect 313 -273 317 -262
rect 329 -269 332 -265
rect 24 -280 347 -273
rect 2 -292 347 -284
rect 2 -360 10 -292
rect 30 -296 35 -292
rect 41 -298 45 -292
rect 65 -298 69 -292
rect 75 -298 79 -292
rect 99 -298 103 -292
rect 109 -298 113 -292
rect 133 -298 137 -292
rect 143 -298 147 -292
rect 167 -298 171 -292
rect 177 -298 181 -292
rect 201 -298 205 -292
rect 211 -298 215 -292
rect 235 -298 239 -292
rect 245 -298 249 -292
rect 269 -298 273 -292
rect 279 -298 283 -292
rect 303 -298 307 -292
rect 313 -298 317 -292
rect 337 -298 341 -292
rect 28 -317 35 -313
rect 53 -314 57 -304
rect 53 -318 65 -314
rect 70 -318 78 -314
rect 87 -315 91 -304
rect 121 -307 125 -304
rect 121 -311 137 -307
rect 28 -325 35 -321
rect 40 -325 44 -321
rect 65 -334 69 -318
rect 87 -319 103 -315
rect 99 -334 103 -319
rect 133 -334 137 -311
rect 155 -314 159 -304
rect 155 -318 171 -314
rect 176 -318 180 -314
rect 189 -317 193 -304
rect 223 -316 227 -304
rect 257 -310 261 -304
rect 291 -308 295 -304
rect 257 -314 282 -310
rect 291 -312 315 -308
rect 167 -334 171 -318
rect 189 -321 205 -317
rect 210 -321 214 -317
rect 223 -320 244 -316
rect 201 -334 205 -321
rect 213 -331 226 -327
rect 235 -334 239 -320
rect 269 -334 273 -314
rect 284 -329 294 -325
rect 303 -334 307 -312
rect 325 -316 329 -304
rect 311 -320 316 -316
rect 325 -320 342 -316
rect 311 -323 315 -320
rect 337 -334 341 -320
rect 41 -349 45 -338
rect 75 -349 79 -338
rect 109 -349 113 -338
rect 143 -349 147 -338
rect 177 -349 181 -338
rect 211 -349 215 -338
rect 245 -349 249 -338
rect 279 -349 283 -338
rect 313 -349 317 -338
rect 329 -345 332 -341
rect 24 -356 347 -349
rect 2 -368 347 -360
rect 2 -436 10 -368
rect 30 -372 35 -368
rect 41 -374 45 -368
rect 65 -374 69 -368
rect 75 -374 79 -368
rect 99 -374 103 -368
rect 109 -374 113 -368
rect 133 -374 137 -368
rect 143 -374 147 -368
rect 167 -374 171 -368
rect 177 -374 181 -368
rect 201 -374 205 -368
rect 211 -374 215 -368
rect 235 -374 239 -368
rect 245 -374 249 -368
rect 269 -374 273 -368
rect 279 -374 283 -368
rect 303 -374 307 -368
rect 313 -374 317 -368
rect 337 -374 341 -368
rect 28 -393 35 -389
rect 53 -390 57 -380
rect 53 -394 65 -390
rect 70 -394 78 -390
rect 87 -391 91 -380
rect 121 -383 125 -380
rect 121 -387 137 -383
rect 28 -401 35 -397
rect 40 -401 44 -397
rect 65 -410 69 -394
rect 87 -395 103 -391
rect 99 -410 103 -395
rect 133 -410 137 -387
rect 155 -390 159 -380
rect 155 -394 171 -390
rect 176 -394 180 -390
rect 189 -393 193 -380
rect 223 -392 227 -380
rect 257 -386 261 -380
rect 291 -384 295 -380
rect 257 -390 282 -386
rect 291 -388 315 -384
rect 167 -410 171 -394
rect 189 -397 205 -393
rect 210 -397 214 -393
rect 223 -396 244 -392
rect 201 -410 205 -397
rect 213 -407 226 -403
rect 235 -410 239 -396
rect 269 -410 273 -390
rect 284 -405 294 -401
rect 303 -410 307 -388
rect 325 -392 329 -380
rect 311 -396 316 -392
rect 325 -396 342 -392
rect 311 -399 315 -396
rect 337 -410 341 -396
rect 41 -425 45 -414
rect 75 -425 79 -414
rect 109 -425 113 -414
rect 143 -425 147 -414
rect 177 -425 181 -414
rect 211 -425 215 -414
rect 245 -425 249 -414
rect 279 -425 283 -414
rect 313 -425 317 -414
rect 329 -421 332 -417
rect 24 -432 347 -425
rect 2 -444 348 -436
rect 2 -511 10 -444
rect 30 -448 35 -444
rect 41 -450 45 -444
rect 65 -450 69 -444
rect 75 -450 79 -444
rect 99 -450 103 -444
rect 109 -450 113 -444
rect 133 -450 137 -444
rect 143 -450 147 -444
rect 167 -450 171 -444
rect 177 -450 181 -444
rect 201 -450 205 -444
rect 211 -450 215 -444
rect 235 -450 239 -444
rect 245 -450 249 -444
rect 269 -450 273 -444
rect 279 -450 283 -444
rect 303 -450 307 -444
rect 313 -450 317 -444
rect 337 -450 341 -444
rect 28 -469 35 -465
rect 53 -466 57 -456
rect 53 -470 65 -466
rect 70 -470 78 -466
rect 87 -467 91 -456
rect 121 -459 125 -456
rect 121 -463 137 -459
rect 28 -477 35 -473
rect 40 -477 44 -473
rect 65 -486 69 -470
rect 87 -471 103 -467
rect 99 -486 103 -471
rect 133 -486 137 -463
rect 155 -466 159 -456
rect 155 -470 171 -466
rect 176 -470 180 -466
rect 189 -469 193 -456
rect 223 -468 227 -456
rect 257 -462 261 -456
rect 291 -460 295 -456
rect 257 -466 282 -462
rect 291 -464 315 -460
rect 167 -486 171 -470
rect 189 -473 205 -469
rect 210 -473 214 -469
rect 223 -472 244 -468
rect 201 -486 205 -473
rect 213 -483 226 -479
rect 235 -486 239 -472
rect 269 -486 273 -466
rect 284 -481 294 -477
rect 303 -486 307 -464
rect 325 -468 329 -456
rect 311 -472 316 -468
rect 325 -472 342 -468
rect 311 -475 315 -472
rect 337 -486 341 -472
rect 41 -501 45 -490
rect 75 -501 79 -490
rect 109 -501 113 -490
rect 143 -501 147 -490
rect 177 -501 181 -490
rect 211 -501 215 -490
rect 245 -501 249 -490
rect 279 -501 283 -490
rect 313 -501 317 -490
rect 329 -497 332 -493
rect 24 -508 347 -501
rect 2 -519 349 -511
rect 2 -520 341 -519
rect 30 -524 35 -520
rect 41 -526 45 -520
rect 65 -526 69 -520
rect 75 -526 79 -520
rect 99 -526 103 -520
rect 109 -526 113 -520
rect 133 -526 137 -520
rect 143 -526 147 -520
rect 167 -526 171 -520
rect 177 -526 181 -520
rect 201 -526 205 -520
rect 211 -526 215 -520
rect 235 -526 239 -520
rect 245 -526 249 -520
rect 269 -526 273 -520
rect 279 -526 283 -520
rect 303 -526 307 -520
rect 313 -526 317 -520
rect 337 -526 341 -520
rect 28 -545 35 -541
rect 53 -542 57 -532
rect 53 -546 65 -542
rect 70 -546 78 -542
rect 87 -543 91 -532
rect 121 -535 125 -532
rect 121 -539 137 -535
rect 28 -553 35 -549
rect 40 -553 44 -549
rect 65 -562 69 -546
rect 87 -547 103 -543
rect 99 -562 103 -547
rect 133 -562 137 -539
rect 155 -542 159 -532
rect 155 -546 171 -542
rect 176 -546 180 -542
rect 189 -545 193 -532
rect 223 -544 227 -532
rect 257 -538 261 -532
rect 291 -536 295 -532
rect 257 -542 282 -538
rect 291 -540 315 -536
rect 167 -562 171 -546
rect 189 -549 205 -545
rect 210 -549 214 -545
rect 223 -548 244 -544
rect 201 -562 205 -549
rect 213 -559 226 -555
rect 235 -562 239 -548
rect 269 -562 273 -542
rect 284 -557 294 -553
rect 303 -562 307 -540
rect 325 -544 329 -532
rect 311 -548 316 -544
rect 325 -548 342 -544
rect 311 -551 315 -548
rect 337 -562 341 -548
rect 41 -577 45 -566
rect 75 -577 79 -566
rect 109 -577 113 -566
rect 143 -577 147 -566
rect 177 -577 181 -566
rect 211 -577 215 -566
rect 245 -577 249 -566
rect 279 -577 283 -566
rect 313 -577 317 -566
rect 329 -573 332 -569
rect -14 -584 347 -577
<< m2contact >>
rect -6 -50 -1 -45
rect 30 8 35 13
rect 35 -13 40 -8
rect 65 -14 70 -9
rect 35 -22 40 -17
rect 51 -22 56 -17
rect 119 -15 124 -10
rect 85 -28 90 -23
rect 103 -26 108 -21
rect 137 -11 142 -6
rect 171 -14 176 -9
rect 243 -8 248 -3
rect 141 -26 146 -21
rect 153 -22 158 -17
rect 205 -17 210 -12
rect 187 -26 192 -21
rect 208 -27 213 -22
rect 244 -17 249 -12
rect 255 -28 260 -23
rect 279 -25 284 -20
rect 342 -16 347 -11
rect 311 -24 316 -19
rect 120 -42 125 -37
rect 324 -42 329 -37
rect 19 -50 24 -45
rect -6 -126 -1 -121
rect 35 -89 40 -84
rect 65 -90 70 -85
rect 35 -98 40 -93
rect 51 -98 56 -93
rect 119 -91 124 -86
rect 85 -104 90 -99
rect 103 -102 108 -97
rect 137 -87 142 -82
rect 171 -90 176 -85
rect 243 -84 248 -79
rect 141 -102 146 -97
rect 153 -98 158 -93
rect 205 -93 210 -88
rect 187 -102 192 -97
rect 208 -103 213 -98
rect 244 -93 249 -88
rect 255 -104 260 -99
rect 279 -101 284 -96
rect 342 -92 347 -87
rect 311 -100 316 -95
rect 120 -118 125 -113
rect 324 -118 329 -113
rect 19 -126 24 -121
rect -6 -202 -1 -197
rect 35 -165 40 -160
rect 65 -166 70 -161
rect 35 -174 40 -169
rect 51 -174 56 -169
rect 119 -167 124 -162
rect 85 -180 90 -175
rect 103 -178 108 -173
rect 137 -163 142 -158
rect 171 -166 176 -161
rect 243 -160 248 -155
rect 141 -178 146 -173
rect 153 -174 158 -169
rect 205 -169 210 -164
rect 187 -178 192 -173
rect 208 -179 213 -174
rect 244 -169 249 -164
rect 255 -180 260 -175
rect 279 -177 284 -172
rect 342 -168 347 -163
rect 311 -176 316 -171
rect 120 -194 125 -189
rect 324 -194 329 -189
rect 19 -202 24 -197
rect -6 -278 -1 -273
rect 35 -241 40 -236
rect 65 -242 70 -237
rect 35 -250 40 -245
rect 51 -250 56 -245
rect 119 -243 124 -238
rect 85 -256 90 -251
rect 103 -254 108 -249
rect 137 -239 142 -234
rect 171 -242 176 -237
rect 243 -236 248 -231
rect 141 -254 146 -249
rect 153 -250 158 -245
rect 205 -245 210 -240
rect 187 -254 192 -249
rect 208 -255 213 -250
rect 244 -245 249 -240
rect 255 -256 260 -251
rect 279 -253 284 -248
rect 342 -244 347 -239
rect 311 -252 316 -247
rect 120 -270 125 -265
rect 324 -270 329 -265
rect 19 -278 24 -273
rect -6 -354 -1 -349
rect 35 -317 40 -312
rect 65 -318 70 -313
rect 35 -326 40 -321
rect 51 -326 56 -321
rect 119 -319 124 -314
rect 85 -332 90 -327
rect 103 -330 108 -325
rect 137 -315 142 -310
rect 171 -318 176 -313
rect 243 -312 248 -307
rect 141 -330 146 -325
rect 153 -326 158 -321
rect 205 -321 210 -316
rect 187 -330 192 -325
rect 208 -331 213 -326
rect 244 -321 249 -316
rect 255 -332 260 -327
rect 279 -329 284 -324
rect 342 -320 347 -315
rect 311 -328 316 -323
rect 120 -346 125 -341
rect 324 -346 329 -341
rect 19 -354 24 -349
rect -6 -430 -1 -425
rect 35 -393 40 -388
rect 65 -394 70 -389
rect 35 -402 40 -397
rect 51 -402 56 -397
rect 119 -395 124 -390
rect 85 -408 90 -403
rect 103 -406 108 -401
rect 137 -391 142 -386
rect 171 -394 176 -389
rect 243 -388 248 -383
rect 141 -406 146 -401
rect 153 -402 158 -397
rect 205 -397 210 -392
rect 187 -406 192 -401
rect 208 -407 213 -402
rect 244 -397 249 -392
rect 255 -408 260 -403
rect 279 -405 284 -400
rect 342 -396 347 -391
rect 311 -404 316 -399
rect 120 -422 125 -417
rect 324 -422 329 -417
rect 19 -430 24 -425
rect -6 -506 -1 -501
rect 35 -469 40 -464
rect 65 -470 70 -465
rect 35 -478 40 -473
rect 51 -478 56 -473
rect 119 -471 124 -466
rect 85 -484 90 -479
rect 103 -482 108 -477
rect 137 -467 142 -462
rect 171 -470 176 -465
rect 243 -464 248 -459
rect 141 -482 146 -477
rect 153 -478 158 -473
rect 205 -473 210 -468
rect 187 -482 192 -477
rect 208 -483 213 -478
rect 244 -473 249 -468
rect 255 -484 260 -479
rect 279 -481 284 -476
rect 342 -472 347 -467
rect 311 -480 316 -475
rect 120 -498 125 -493
rect 324 -498 329 -493
rect 19 -506 24 -501
rect 35 -545 40 -540
rect 65 -546 70 -541
rect 35 -554 40 -549
rect 51 -554 56 -549
rect 119 -547 124 -542
rect 85 -560 90 -555
rect 103 -558 108 -553
rect 137 -543 142 -538
rect 171 -546 176 -541
rect 243 -540 248 -535
rect 141 -558 146 -553
rect 153 -554 158 -549
rect 205 -549 210 -544
rect 187 -558 192 -553
rect 208 -559 213 -554
rect 244 -549 249 -544
rect 255 -560 260 -555
rect 279 -557 284 -552
rect 342 -548 347 -543
rect 311 -556 316 -551
rect 120 -574 125 -569
rect 324 -574 329 -569
<< metal2 >>
rect 35 9 243 13
rect 36 -5 109 -1
rect 36 -8 40 -5
rect 40 -13 55 -9
rect 51 -17 55 -13
rect 105 -10 109 -5
rect 105 -14 119 -10
rect 66 -15 70 -14
rect 142 -11 158 -7
rect 66 -19 99 -15
rect 154 -17 158 -11
rect 36 -38 40 -22
rect 70 -28 85 -24
rect 70 -38 74 -28
rect 36 -42 74 -38
rect 95 -42 99 -19
rect 108 -26 141 -22
rect 172 -30 176 -14
rect 187 -21 191 9
rect 206 -8 227 -4
rect 239 -8 243 9
rect 206 -12 210 -8
rect 223 -17 227 -8
rect 249 -17 283 -13
rect 223 -21 239 -17
rect 235 -23 239 -21
rect 279 -20 283 -17
rect 235 -27 255 -23
rect 208 -30 212 -27
rect 172 -34 212 -30
rect 255 -30 260 -28
rect 311 -30 315 -24
rect 255 -34 315 -30
rect -1 -50 19 -45
rect 95 -46 329 -42
rect 343 -64 347 -16
rect 187 -69 347 -64
rect 36 -81 109 -77
rect 36 -84 40 -81
rect 40 -89 55 -85
rect 51 -93 55 -89
rect 105 -86 109 -81
rect 105 -90 119 -86
rect 66 -91 70 -90
rect 142 -87 158 -83
rect 66 -95 99 -91
rect 154 -93 158 -87
rect 36 -114 40 -98
rect 70 -104 85 -100
rect 70 -114 74 -104
rect 36 -118 74 -114
rect 95 -118 99 -95
rect 108 -102 141 -98
rect 172 -106 176 -90
rect 187 -97 191 -69
rect 206 -84 227 -80
rect 239 -84 243 -69
rect 206 -88 210 -84
rect 223 -93 227 -84
rect 249 -93 283 -89
rect 223 -97 239 -93
rect 235 -99 239 -97
rect 279 -96 283 -93
rect 235 -103 255 -99
rect 208 -106 212 -103
rect 172 -110 212 -106
rect 255 -106 260 -104
rect 311 -106 315 -100
rect 255 -110 315 -106
rect -1 -126 19 -121
rect 95 -122 329 -118
rect 342 -143 347 -92
rect 186 -148 347 -143
rect 36 -157 109 -153
rect 36 -160 40 -157
rect 40 -165 55 -161
rect 51 -169 55 -165
rect 105 -162 109 -157
rect 105 -166 119 -162
rect 66 -167 70 -166
rect 142 -163 158 -159
rect 66 -171 99 -167
rect 154 -169 158 -163
rect 36 -190 40 -174
rect 70 -180 85 -176
rect 70 -190 74 -180
rect 36 -194 74 -190
rect 95 -194 99 -171
rect 108 -178 141 -174
rect 172 -182 176 -166
rect 187 -173 191 -148
rect 206 -160 227 -156
rect 239 -160 243 -148
rect 342 -149 347 -148
rect 206 -164 210 -160
rect 223 -169 227 -160
rect 249 -169 283 -165
rect 223 -173 239 -169
rect 235 -175 239 -173
rect 279 -172 283 -169
rect 235 -179 255 -175
rect 208 -182 212 -179
rect 172 -186 212 -182
rect 255 -182 260 -180
rect 311 -182 315 -176
rect 255 -186 315 -182
rect -1 -202 19 -197
rect 95 -198 329 -194
rect 342 -220 347 -168
rect 186 -225 347 -220
rect 36 -233 109 -229
rect 36 -236 40 -233
rect 40 -241 55 -237
rect 51 -245 55 -241
rect 105 -238 109 -233
rect 105 -242 119 -238
rect 66 -243 70 -242
rect 142 -239 158 -235
rect 66 -247 99 -243
rect 154 -245 158 -239
rect 36 -266 40 -250
rect 70 -256 85 -252
rect 70 -266 74 -256
rect 36 -270 74 -266
rect 95 -270 99 -247
rect 108 -254 141 -250
rect 172 -258 176 -242
rect 187 -249 191 -225
rect 206 -236 227 -232
rect 239 -236 243 -225
rect 206 -240 210 -236
rect 223 -245 227 -236
rect 249 -245 283 -241
rect 223 -249 239 -245
rect 235 -251 239 -249
rect 279 -248 283 -245
rect 235 -255 255 -251
rect 208 -258 212 -255
rect 172 -262 212 -258
rect 255 -258 260 -256
rect 311 -258 315 -252
rect 255 -262 315 -258
rect -1 -278 19 -273
rect 95 -274 329 -270
rect 342 -296 347 -244
rect 187 -301 347 -296
rect 36 -309 109 -305
rect 36 -312 40 -309
rect 40 -317 55 -313
rect 51 -321 55 -317
rect 105 -314 109 -309
rect 105 -318 119 -314
rect 66 -319 70 -318
rect 142 -315 158 -311
rect 66 -323 99 -319
rect 154 -321 158 -315
rect 36 -342 40 -326
rect 70 -332 85 -328
rect 70 -342 74 -332
rect 36 -346 74 -342
rect 95 -346 99 -323
rect 108 -330 141 -326
rect 172 -334 176 -318
rect 187 -325 191 -301
rect 206 -312 227 -308
rect 239 -312 243 -301
rect 206 -316 210 -312
rect 223 -321 227 -312
rect 249 -321 283 -317
rect 223 -325 239 -321
rect 235 -327 239 -325
rect 279 -324 283 -321
rect 235 -331 255 -327
rect 208 -334 212 -331
rect 172 -338 212 -334
rect 255 -334 260 -332
rect 311 -334 315 -328
rect 255 -338 315 -334
rect -1 -354 19 -349
rect 95 -350 329 -346
rect 342 -373 347 -320
rect 186 -378 347 -373
rect 36 -385 109 -381
rect 36 -388 40 -385
rect 40 -393 55 -389
rect 51 -397 55 -393
rect 105 -390 109 -385
rect 105 -394 119 -390
rect 66 -395 70 -394
rect 142 -391 158 -387
rect 66 -399 99 -395
rect 154 -397 158 -391
rect 36 -418 40 -402
rect 70 -408 85 -404
rect 70 -418 74 -408
rect 36 -422 74 -418
rect 95 -422 99 -399
rect 108 -406 141 -402
rect 172 -410 176 -394
rect 187 -401 191 -378
rect 206 -388 227 -384
rect 239 -388 243 -378
rect 206 -392 210 -388
rect 223 -397 227 -388
rect 249 -397 283 -393
rect 223 -401 239 -397
rect 235 -403 239 -401
rect 279 -400 283 -397
rect 235 -407 255 -403
rect 208 -410 212 -407
rect 172 -414 212 -410
rect 255 -410 260 -408
rect 311 -410 315 -404
rect 255 -414 315 -410
rect -1 -430 19 -425
rect 95 -426 329 -422
rect 342 -448 347 -396
rect 186 -453 347 -448
rect 36 -461 109 -457
rect 36 -464 40 -461
rect 40 -469 55 -465
rect 51 -473 55 -469
rect 105 -466 109 -461
rect 105 -470 119 -466
rect 66 -471 70 -470
rect 142 -467 158 -463
rect 66 -475 99 -471
rect 154 -473 158 -467
rect 36 -494 40 -478
rect 70 -484 85 -480
rect 70 -494 74 -484
rect 36 -498 74 -494
rect 95 -498 99 -475
rect 108 -482 141 -478
rect 172 -486 176 -470
rect 187 -477 191 -453
rect 206 -464 227 -460
rect 239 -464 243 -453
rect 206 -468 210 -464
rect 223 -473 227 -464
rect 249 -473 283 -469
rect 223 -477 239 -473
rect 235 -479 239 -477
rect 279 -476 283 -473
rect 235 -483 255 -479
rect 208 -486 212 -483
rect 172 -490 212 -486
rect 255 -486 260 -484
rect 311 -486 315 -480
rect 255 -490 315 -486
rect -1 -506 19 -501
rect 95 -502 329 -498
rect 342 -523 347 -472
rect 186 -528 347 -523
rect 36 -537 109 -533
rect 36 -540 40 -537
rect 40 -545 55 -541
rect 51 -549 55 -545
rect 105 -542 109 -537
rect 105 -546 119 -542
rect 66 -547 70 -546
rect 142 -543 158 -539
rect 66 -551 99 -547
rect 154 -549 158 -543
rect 36 -570 40 -554
rect 70 -560 85 -556
rect 70 -570 74 -560
rect 36 -574 74 -570
rect 95 -574 99 -551
rect 108 -558 141 -554
rect 172 -562 176 -546
rect 187 -553 191 -528
rect 206 -540 227 -536
rect 239 -540 243 -528
rect 206 -544 210 -540
rect 223 -549 227 -540
rect 249 -549 283 -545
rect 223 -553 239 -549
rect 235 -555 239 -553
rect 279 -552 283 -549
rect 235 -559 255 -555
rect 208 -562 212 -559
rect 172 -566 212 -562
rect 255 -562 260 -560
rect 311 -562 315 -556
rect 255 -566 315 -562
rect 95 -578 329 -574
<< labels >>
rlabel metal1 6 18 6 18 4 Vdd
rlabel metal1 -10 18 -10 18 3 Gnd
rlabel metal1 31 -11 31 -11 1 b0
rlabel metal1 30 -19 30 -19 1 a0
rlabel metal1 30 6 30 6 1 cin0
rlabel metal1 312 -6 312 -6 1 sum0
rlabel metal1 31 -87 31 -87 1 b1
rlabel metal1 31 -95 31 -95 1 a1
rlabel metal1 312 -82 312 -82 1 sum1
rlabel metal1 306 -159 306 -159 1 sum2
rlabel metal1 30 -162 30 -162 1 b2
rlabel metal1 29 -171 29 -171 1 a2
rlabel metal1 31 -239 31 -239 1 b3
rlabel metal1 30 -248 30 -248 1 a3
rlabel metal1 309 -234 309 -234 1 sum3
rlabel metal1 29 -316 29 -316 1 b4
rlabel metal1 30 -324 30 -324 1 a4
rlabel metal1 312 -310 312 -310 1 sum4
rlabel metal1 30 -391 30 -391 1 b5
rlabel metal1 29 -399 29 -399 1 a5
rlabel metal1 310 -386 310 -386 1 sum5
rlabel metal1 30 -467 30 -467 1 b6
rlabel metal1 32 -476 32 -476 1 a6
rlabel metal1 312 -462 312 -462 1 sum6
rlabel metal1 31 -543 31 -543 1 b7
rlabel metal1 30 -552 30 -552 1 a7
rlabel metal1 312 -537 312 -537 1 sum7
rlabel metal1 340 -545 340 -545 1 cout7
<< end >>
